library ieee;
use ieee.std_logic_1164.all;

entity partial_products_add is
	--port();
end entity;

architecture beh of partial_products_add is
begin

end architecture;
