library ieee;
use ieee.std_logic_1164.all;
use work.pp_array_pkg.all;


entity daddaTree is
        port(   pp_ext: in ppmatrix;
                        Addend1: out std_logic_vector(63 downto 0);
                        Addend2: out std_logic_vector(63 downto 0));
end entity;

architecture rtl of daddaTree is
        component full_adder is
                port(   A,B,Cin: in std_logic;
                        S,Cout: out std_logic);
        end component full_adder;
        component half_adder is
                port(   A,B: in std_logic;
                        S,Cout: out std_logic);
        end component half_adder;


signal resultHA0, carryOutHA0, resultHA1, carryOutHA1, resultFA0, carryOutFA0, resultHA2, carryOutHA2, resultFA1, carryOutFA1, resultHA3, carryOutHA3, resultFA2, carryOutFA2, resultFA3, carryOutFA3, resultHA4, carryOutHA4, resultFA4, carryOutFA4, resultFA5, carryOutFA5, resultHA5, carryOutHA5, resultFA6, carryOutFA6, resultFA7, carryOutFA7, resultFA8, carryOutFA8, resultHA6, carryOutHA6, resultFA9, carryOutFA9, resultFA10, carryOutFA10, resultFA11, carryOutFA11, resultHA7, carryOutHA7, resultFA12, carryOutFA12, resultFA13, carryOutFA13, resultFA14, carryOutFA14, resultFA15, carryOutFA15, resultFA16, carryOutFA16, resultFA17, carryOutFA17, resultFA18, carryOutFA18, resultFA19, carryOutFA19, resultFA20, carryOutFA20, resultFA21, carryOutFA21, resultFA22, carryOutFA22, resultFA23, carryOutFA23, resultFA24, carryOutFA24, resultFA25, carryOutFA25, resultFA26, carryOutFA26, resultFA27, carryOutFA27, resultFA28, carryOutFA28, resultFA29, carryOutFA29, resultFA30, carryOutFA30, resultHA8, carryOutHA8, resultFA31, carryOutFA31, resultFA32, carryOutFA32, resultFA33, carryOutFA33, resultFA34, carryOutFA34, resultFA35, carryOutFA35, resultHA9, carryOutHA9, resultFA36, carryOutFA36, resultFA37, carryOutFA37, resultFA38, carryOutFA38, resultHA10, carryOutHA10, resultFA39, carryOutFA39, resultHA11, carryOutHA11, resultHA12, carryOutHA12, resultHA13, carryOutHA13, resultFA40, carryOutFA40, resultHA14, carryOutHA14, resultFA41, carryOutFA41, resultHA15, carryOutHA15, resultFA42, carryOutFA42, resultFA43, carryOutFA43, resultHA16, carryOutHA16, resultFA44, carryOutFA44, resultFA45, carryOutFA45, resultHA17, carryOutHA17, resultFA46, carryOutFA46, resultFA47, carryOutFA47, resultFA48, carryOutFA48, resultHA18, carryOutHA18, resultFA49, carryOutFA49, resultFA50, carryOutFA50, resultFA51, carryOutFA51, resultHA19, carryOutHA19, resultFA52, carryOutFA52, resultFA53, carryOutFA53, resultFA54, carryOutFA54, resultFA55, carryOutFA55, resultFA56, carryOutFA56, resultFA57, carryOutFA57, resultFA58, carryOutFA58, resultFA59, carryOutFA59, resultFA60, carryOutFA60, resultFA61, carryOutFA61, resultFA62, carryOutFA62, resultFA63, carryOutFA63, resultFA64, carryOutFA64, resultFA65, carryOutFA65, resultFA66, carryOutFA66, resultFA67, carryOutFA67, resultFA68, carryOutFA68, resultFA69, carryOutFA69, resultFA70, carryOutFA70, resultFA71, carryOutFA71, resultFA72, carryOutFA72, resultFA73, carryOutFA73, resultFA74, carryOutFA74, resultFA75, carryOutFA75, resultFA76, carryOutFA76, resultFA77, carryOutFA77, resultFA78, carryOutFA78, resultFA79, carryOutFA79, resultFA80, carryOutFA80, resultFA81, carryOutFA81, resultFA82, carryOutFA82, resultFA83, carryOutFA83, resultFA84, carryOutFA84, resultFA85, carryOutFA85, resultFA86, carryOutFA86, resultFA87, carryOutFA87, resultFA88, carryOutFA88, resultFA89, carryOutFA89, resultFA90, carryOutFA90, resultFA91, carryOutFA91, resultFA92, carryOutFA92, resultFA93, carryOutFA93, resultFA94, carryOutFA94, resultFA95, carryOutFA95, resultFA96, carryOutFA96, resultFA97, carryOutFA97, resultFA98, carryOutFA98, resultFA99, carryOutFA99, resultFA100, carryOutFA100, resultFA101, carryOutFA101, resultFA102, carryOutFA102, resultFA103, carryOutFA103, resultFA104, carryOutFA104, resultFA105, carryOutFA105, resultFA106, carryOutFA106, resultFA107, carryOutFA107, resultFA108, carryOutFA108, resultFA109, carryOutFA109, resultFA110, carryOutFA110, resultFA111, carryOutFA111, resultFA112, carryOutFA112, resultFA113, carryOutFA113, resultFA114, carryOutFA114, resultFA115, carryOutFA115, resultFA116, carryOutFA116, resultFA117, carryOutFA117, resultFA118, carryOutFA118, resultFA119, carryOutFA119, resultFA120, carryOutFA120, resultFA121, carryOutFA121, resultFA122, carryOutFA122, resultFA123, carryOutFA123, resultFA124, carryOutFA124, resultFA125, carryOutFA125, resultFA126, carryOutFA126, resultFA127, carryOutFA127, resultFA128, carryOutFA128, resultFA129, carryOutFA129, resultFA130, carryOutFA130, resultFA131, carryOutFA131, resultFA132, carryOutFA132, resultFA133, carryOutFA133, resultFA134, carryOutFA134, resultHA20, carryOutHA20, resultFA135, carryOutFA135, resultFA136, carryOutFA136, resultFA137, carryOutFA137, resultFA138, carryOutFA138, resultFA139, carryOutFA139, resultHA21, carryOutHA21, resultFA140, carryOutFA140, resultFA141, carryOutFA141, resultFA142, carryOutFA142, resultHA22, carryOutHA22, resultFA143, carryOutFA143, resultHA23, carryOutHA23, resultHA24, carryOutHA24, resultHA25, carryOutHA25, resultFA144, carryOutFA144, resultHA26, carryOutHA26, resultFA145, carryOutFA145, resultHA27, carryOutHA27, resultFA146, carryOutFA146, resultFA147, carryOutFA147, resultHA28, carryOutHA28, resultFA148, carryOutFA148, resultFA149, carryOutFA149, resultHA29, carryOutHA29, resultFA150, carryOutFA150, resultFA151, carryOutFA151, resultFA152, carryOutFA152, resultFA153, carryOutFA153, resultFA154, carryOutFA154, resultFA155, carryOutFA155, resultFA156, carryOutFA156, resultFA157, carryOutFA157, resultFA158, carryOutFA158, resultFA159, carryOutFA159, resultFA160, carryOutFA160, resultFA161, carryOutFA161, resultFA162, carryOutFA162, resultFA163, carryOutFA163, resultFA164, carryOutFA164, resultFA165, carryOutFA165, resultFA166, carryOutFA166, resultFA167, carryOutFA167, resultFA168, carryOutFA168, resultFA169, carryOutFA169, resultFA170, carryOutFA170, resultFA171, carryOutFA171, resultFA172, carryOutFA172, resultFA173, carryOutFA173, resultFA174, carryOutFA174, resultFA175, carryOutFA175, resultFA176, carryOutFA176, resultFA177, carryOutFA177, resultFA178, carryOutFA178, resultFA179, carryOutFA179, resultFA180, carryOutFA180, resultFA181, carryOutFA181, resultFA182, carryOutFA182, resultFA183, carryOutFA183, resultFA184, carryOutFA184, resultFA185, carryOutFA185, resultFA186, carryOutFA186, resultFA187, carryOutFA187, resultFA188, carryOutFA188, resultFA189, carryOutFA189, resultFA190, carryOutFA190, resultFA191, carryOutFA191, resultFA192, carryOutFA192, resultFA193, carryOutFA193, resultFA194, carryOutFA194, resultFA195, carryOutFA195, resultFA196, carryOutFA196, resultFA197, carryOutFA197, resultFA198, carryOutFA198, resultFA199, carryOutFA199, resultFA200, carryOutFA200, resultFA201, carryOutFA201, resultFA202, carryOutFA202, resultFA203, carryOutFA203, resultFA204, carryOutFA204, resultFA205, carryOutFA205, resultFA206, carryOutFA206, resultFA207, carryOutFA207, resultFA208, carryOutFA208, resultFA209, carryOutFA209, resultFA210, carryOutFA210, resultFA211, carryOutFA211, resultFA212, carryOutFA212, resultFA213, carryOutFA213, resultFA214, carryOutFA214, resultFA215, carryOutFA215, resultFA216, carryOutFA216, resultFA217, carryOutFA217, resultFA218, carryOutFA218, resultFA219, carryOutFA219, resultFA220, carryOutFA220, resultFA221, carryOutFA221, resultFA222, carryOutFA222, resultFA223, carryOutFA223, resultFA224, carryOutFA224, resultFA225, carryOutFA225, resultFA226, carryOutFA226, resultFA227, carryOutFA227, resultFA228, carryOutFA228, resultFA229, carryOutFA229, resultFA230, carryOutFA230, resultFA231, carryOutFA231, resultFA232, carryOutFA232, resultFA233, carryOutFA233, resultFA234, carryOutFA234, resultFA235, carryOutFA235, resultFA236, carryOutFA236, resultFA237, carryOutFA237, resultFA238, carryOutFA238, resultFA239, carryOutFA239, resultFA240, carryOutFA240, resultFA241, carryOutFA241, resultFA242, carryOutFA242, resultFA243, carryOutFA243, resultFA244, carryOutFA244, resultFA245, carryOutFA245, resultFA246, carryOutFA246, resultFA247, carryOutFA247, resultFA248, carryOutFA248, resultFA249, carryOutFA249, resultFA250, carryOutFA250, resultFA251, carryOutFA251, resultFA252, carryOutFA252, resultFA253, carryOutFA253, resultFA254, carryOutFA254, resultFA255, carryOutFA255, resultFA256, carryOutFA256, resultFA257, carryOutFA257, resultFA258, carryOutFA258, resultFA259, carryOutFA259, resultHA30, carryOutHA30, resultFA260, carryOutFA260, resultFA261, carryOutFA261, resultFA262, carryOutFA262, resultHA31, carryOutHA31, resultFA263, carryOutFA263, resultHA32, carryOutHA32, resultHA33, carryOutHA33, resultHA34, carryOutHA34, resultFA264, carryOutFA264, resultHA35, carryOutHA35, resultFA265, carryOutFA265, resultHA36, carryOutHA36, resultFA266, carryOutFA266, resultFA267, carryOutFA267, resultFA268, carryOutFA268, resultFA269, carryOutFA269, resultFA270, carryOutFA270, resultFA271, carryOutFA271, resultFA272, carryOutFA272, resultFA273, carryOutFA273, resultFA274, carryOutFA274, resultFA275, carryOutFA275, resultFA276, carryOutFA276, resultFA277, carryOutFA277, resultFA278, carryOutFA278, resultFA279, carryOutFA279, resultFA280, carryOutFA280, resultFA281, carryOutFA281, resultFA282, carryOutFA282, resultFA283, carryOutFA283, resultFA284, carryOutFA284, resultFA285, carryOutFA285, resultFA286, carryOutFA286, resultFA287, carryOutFA287, resultFA288, carryOutFA288, resultFA289, carryOutFA289, resultFA290, carryOutFA290, resultFA291, carryOutFA291, resultFA292, carryOutFA292, resultFA293, carryOutFA293, resultFA294, carryOutFA294, resultFA295, carryOutFA295, resultFA296, carryOutFA296, resultFA297, carryOutFA297, resultFA298, carryOutFA298, resultFA299, carryOutFA299, resultFA300, carryOutFA300, resultFA301, carryOutFA301, resultFA302, carryOutFA302, resultFA303, carryOutFA303, resultFA304, carryOutFA304, resultFA305, carryOutFA305, resultFA306, carryOutFA306, resultFA307, carryOutFA307, resultFA308, carryOutFA308, resultFA309, carryOutFA309, resultFA310, carryOutFA310, resultFA311, carryOutFA311, resultFA312, carryOutFA312, resultFA313, carryOutFA313, resultFA314, carryOutFA314, resultFA315, carryOutFA315, resultFA316, carryOutFA316, resultFA317, carryOutFA317, resultFA318, carryOutFA318, resultFA319, carryOutFA319, resultFA320, carryOutFA320, resultFA321, carryOutFA321, resultFA322, carryOutFA322, resultFA323, carryOutFA323, resultFA324, carryOutFA324, resultFA325, carryOutFA325, resultFA326, carryOutFA326, resultFA327, carryOutFA327, resultFA328, carryOutFA328, resultFA329, carryOutFA329, resultFA330, carryOutFA330, resultFA331, carryOutFA331, resultFA332, carryOutFA332, resultFA333, carryOutFA333, resultFA334, carryOutFA334, resultFA335, carryOutFA335, resultFA336, carryOutFA336, resultFA337, carryOutFA337, resultFA338, carryOutFA338, resultFA339, carryOutFA339, resultFA340, carryOutFA340, resultFA341, carryOutFA341, resultFA342, carryOutFA342, resultFA343, carryOutFA343, resultFA344, carryOutFA344, resultFA345, carryOutFA345, resultFA346, carryOutFA346, resultFA347, carryOutFA347, resultFA348, carryOutFA348, resultFA349, carryOutFA349, resultFA350, carryOutFA350, resultFA351, carryOutFA351, resultFA352, carryOutFA352, resultFA353, carryOutFA353, resultFA354, carryOutFA354, resultFA355, carryOutFA355, resultFA356, carryOutFA356, resultFA357, carryOutFA357, resultFA358, carryOutFA358, resultFA359, carryOutFA359, resultFA360, carryOutFA360, resultFA361, carryOutFA361, resultFA362, carryOutFA362, resultHA37, carryOutHA37, resultFA363, carryOutFA363, resultHA38, carryOutHA38, resultHA39, carryOutHA39, resultHA40, carryOutHA40, resultFA364, carryOutFA364, resultFA365, carryOutFA365, resultFA366, carryOutFA366, resultFA367, carryOutFA367, resultFA368, carryOutFA368, resultFA369, carryOutFA369, resultFA370, carryOutFA370, resultFA371, carryOutFA371, resultFA372, carryOutFA372, resultFA373, carryOutFA373, resultFA374, carryOutFA374, resultFA375, carryOutFA375, resultFA376, carryOutFA376, resultFA377, carryOutFA377, resultFA378, carryOutFA378, resultFA379, carryOutFA379, resultFA380, carryOutFA380, resultFA381, carryOutFA381, resultFA382, carryOutFA382, resultFA383, carryOutFA383, resultFA384, carryOutFA384, resultFA385, carryOutFA385, resultFA386, carryOutFA386, resultFA387, carryOutFA387, resultFA388, carryOutFA388, resultFA389, carryOutFA389, resultFA390, carryOutFA390, resultFA391, carryOutFA391, resultFA392, carryOutFA392, resultFA393, carryOutFA393, resultFA394, carryOutFA394, resultFA395, carryOutFA395, resultFA396, carryOutFA396, resultFA397, carryOutFA397, resultFA398, carryOutFA398, resultFA399, carryOutFA399, resultFA400, carryOutFA400, resultFA401, carryOutFA401, resultFA402, carryOutFA402, resultFA403, carryOutFA403, resultFA404, carryOutFA404, resultFA405, carryOutFA405, resultFA406, carryOutFA406, resultFA407, carryOutFA407, resultFA408, carryOutFA408, resultFA409, carryOutFA409, resultFA410, carryOutFA410, resultFA411, carryOutFA411, resultFA412, carryOutFA412, resultFA413, carryOutFA413, resultFA414, carryOutFA414, resultFA415, carryOutFA415, resultFA416, carryOutFA416, resultFA417, carryOutFA417, resultFA418, carryOutFA418, resultFA419, carryOutFA419, resultHA41, carryOutHA41, resultHA42, carryOutHA42, resultHA43, carryOutHA43, resultFA420, carryOutFA420, resultFA421, carryOutFA421, resultFA422, carryOutFA422, resultFA423, carryOutFA423, resultFA424, carryOutFA424, resultFA425, carryOutFA425, resultFA426, carryOutFA426, resultFA427, carryOutFA427, resultFA428, carryOutFA428, resultFA429, carryOutFA429, resultFA430, carryOutFA430, resultFA431, carryOutFA431, resultFA432, carryOutFA432, resultFA433, carryOutFA433, resultFA434, carryOutFA434, resultFA435, carryOutFA435, resultFA436, carryOutFA436, resultFA437, carryOutFA437, resultFA438, carryOutFA438, resultFA439, carryOutFA439, resultFA440, carryOutFA440, resultFA441, carryOutFA441, resultFA442, carryOutFA442, resultFA443, carryOutFA443, resultFA444, carryOutFA444, resultFA445, carryOutFA445, resultFA446, carryOutFA446, resultFA447, carryOutFA447, resultFA448, carryOutFA448, resultFA449, carryOutFA449, resultFA450, carryOutFA450, resultFA451, carryOutFA451, resultFA452, carryOutFA452, resultFA453, carryOutFA453, resultFA454, carryOutFA454, resultFA455, carryOutFA455, resultFA456, carryOutFA456, resultFA457, carryOutFA457, resultFA458, carryOutFA458, resultFA459, carryOutFA459, resultFA460, carryOutFA460, resultFA461, carryOutFA461, resultFA462, carryOutFA462, resultFA463, carryOutFA463, resultFA464, carryOutFA464, resultFA465, carryOutFA465, resultFA466, carryOutFA466, resultFA467, carryOutFA467, resultFA468, carryOutFA468, resultFA469, carryOutFA469, resultFA470, carryOutFA470, resultFA471, carryOutFA471, resultFA472, carryOutFA472, resultFA473, carryOutFA473, resultFA474, carryOutFA474, resultFA475, carryOutFA475, resultFA476, carryOutFA476, resultFA477, carryOutFA477, resultFA478, carryOutFA478, resultFA479, carryOutFA479: std_logic;
begin
HA0:half_adder port map (A => pp_ext(0)(24), B => pp_ext(1)(24), S => resultHA0, Cout => carryOutHA0);
HA1:half_adder port map (A => pp_ext(0)(25), B => pp_ext(1)(25), S => resultHA1, Cout => carryOutHA1);
FA0:full_adder port map (A => pp_ext(0)(26), B => pp_ext(1)(26), Cin => pp_ext(2)(24), S => resultFA0, Cout => carryOutFA0);
HA2:half_adder port map (A => pp_ext(3)(22), B => pp_ext(4)(20), S => resultHA2, Cout => carryOutHA2);
FA1:full_adder port map (A => pp_ext(0)(27), B => pp_ext(1)(27), Cin => pp_ext(2)(25), S => resultFA1, Cout => carryOutFA1);
HA3:half_adder port map (A => pp_ext(3)(23), B => pp_ext(4)(21), S => resultHA3, Cout => carryOutHA3);
FA2:full_adder port map (A => pp_ext(0)(28), B => pp_ext(1)(28), Cin => pp_ext(2)(26), S => resultFA2, Cout => carryOutFA2);
FA3:full_adder port map (A => pp_ext(3)(24), B => pp_ext(4)(22), Cin => pp_ext(5)(20), S => resultFA3, Cout => carryOutFA3);
HA4:half_adder port map (A => pp_ext(6)(18), B => pp_ext(7)(16), S => resultHA4, Cout => carryOutHA4);
FA4:full_adder port map (A => pp_ext(0)(29), B => pp_ext(1)(29), Cin => pp_ext(2)(27), S => resultFA4, Cout => carryOutFA4);
FA5:full_adder port map (A => pp_ext(3)(25), B => pp_ext(4)(23), Cin => pp_ext(5)(21), S => resultFA5, Cout => carryOutFA5);
HA5:half_adder port map (A => pp_ext(6)(19), B => pp_ext(7)(17), S => resultHA5, Cout => carryOutHA5);
FA6:full_adder port map (A => pp_ext(0)(30), B => pp_ext(1)(30), Cin => pp_ext(2)(28), S => resultFA6, Cout => carryOutFA6);
FA7:full_adder port map (A => pp_ext(3)(26), B => pp_ext(4)(24), Cin => pp_ext(5)(22), S => resultFA7, Cout => carryOutFA7);
FA8:full_adder port map (A => pp_ext(6)(20), B => pp_ext(7)(18), Cin => pp_ext(8)(16), S => resultFA8, Cout => carryOutFA8);
HA6:half_adder port map (A => pp_ext(9)(14), B => pp_ext(10)(12), S => resultHA6, Cout => carryOutHA6);
FA9:full_adder port map (A => pp_ext(0)(31), B => pp_ext(1)(31), Cin => pp_ext(2)(29), S => resultFA9, Cout => carryOutFA9);
FA10:full_adder port map (A => pp_ext(3)(27), B => pp_ext(4)(25), Cin => pp_ext(5)(23), S => resultFA10, Cout => carryOutFA10);
FA11:full_adder port map (A => pp_ext(6)(21), B => pp_ext(7)(19), Cin => pp_ext(8)(17), S => resultFA11, Cout => carryOutFA11);
HA7:half_adder port map (A => pp_ext(9)(15), B => pp_ext(10)(13), S => resultHA7, Cout => carryOutHA7);
FA12:full_adder port map (A => pp_ext(0)(32), B => pp_ext(1)(32), Cin => pp_ext(2)(30), S => resultFA12, Cout => carryOutFA12);
FA13:full_adder port map (A => pp_ext(3)(28), B => pp_ext(4)(26), Cin => pp_ext(5)(24), S => resultFA13, Cout => carryOutFA13);
FA14:full_adder port map (A => pp_ext(6)(22), B => pp_ext(7)(20), Cin => pp_ext(8)(18), S => resultFA14, Cout => carryOutFA14);
FA15:full_adder port map (A => pp_ext(9)(16), B => pp_ext(10)(14), Cin => pp_ext(11)(12), S => resultFA15, Cout => carryOutFA15);
FA16:full_adder port map (A => pp_ext(0)(33), B => pp_ext(1)(33), Cin => pp_ext(2)(31), S => resultFA16, Cout => carryOutFA16);
FA17:full_adder port map (A => pp_ext(3)(29), B => pp_ext(4)(27), Cin => pp_ext(5)(25), S => resultFA17, Cout => carryOutFA17);
FA18:full_adder port map (A => pp_ext(6)(23), B => pp_ext(7)(21), Cin => pp_ext(8)(19), S => resultFA18, Cout => carryOutFA18);
FA19:full_adder port map (A => pp_ext(9)(17), B => pp_ext(10)(15), Cin => pp_ext(11)(13), S => resultFA19, Cout => carryOutFA19);
FA20:full_adder port map (A => pp_ext(0)(34), B => pp_ext(1)(34), Cin => pp_ext(2)(32), S => resultFA20, Cout => carryOutFA20);
FA21:full_adder port map (A => pp_ext(3)(30), B => pp_ext(4)(28), Cin => pp_ext(5)(26), S => resultFA21, Cout => carryOutFA21);
FA22:full_adder port map (A => pp_ext(6)(24), B => pp_ext(7)(22), Cin => pp_ext(8)(20), S => resultFA22, Cout => carryOutFA22);
FA23:full_adder port map (A => pp_ext(9)(18), B => pp_ext(10)(16), Cin => pp_ext(11)(14), S => resultFA23, Cout => carryOutFA23);
FA24:full_adder port map (A => pp_ext(0)(35), B => pp_ext(1)(35), Cin => pp_ext(2)(33), S => resultFA24, Cout => carryOutFA24);
FA25:full_adder port map (A => pp_ext(3)(31), B => pp_ext(4)(29), Cin => pp_ext(5)(27), S => resultFA25, Cout => carryOutFA25);
FA26:full_adder port map (A => pp_ext(6)(25), B => pp_ext(7)(23), Cin => pp_ext(8)(21), S => resultFA26, Cout => carryOutFA26);
FA27:full_adder port map (A => pp_ext(9)(19), B => pp_ext(10)(17), Cin => pp_ext(11)(15), S => resultFA27, Cout => carryOutFA27);
FA28:full_adder port map (A => pp_ext(1)(36), B => pp_ext(2)(34), Cin => pp_ext(3)(32), S => resultFA28, Cout => carryOutFA28);
FA29:full_adder port map (A => pp_ext(4)(30), B => pp_ext(5)(28), Cin => pp_ext(6)(26), S => resultFA29, Cout => carryOutFA29);
FA30:full_adder port map (A => pp_ext(7)(24), B => pp_ext(8)(22), Cin => pp_ext(9)(20), S => resultFA30, Cout => carryOutFA30);
HA8:half_adder port map (A => pp_ext(10)(18), B => pp_ext(11)(16), S => resultHA8, Cout => carryOutHA8);
FA31:full_adder port map (A => pp_ext(2)(35), B => pp_ext(3)(33), Cin => pp_ext(4)(31), S => resultFA31, Cout => carryOutFA31);
FA32:full_adder port map (A => pp_ext(5)(29), B => pp_ext(6)(27), Cin => pp_ext(7)(25), S => resultFA32, Cout => carryOutFA32);
FA33:full_adder port map (A => pp_ext(8)(23), B => pp_ext(9)(21), Cin => pp_ext(10)(19), S => resultFA33, Cout => carryOutFA33);
FA34:full_adder port map (A => pp_ext(2)(36), B => pp_ext(3)(34), Cin => pp_ext(4)(32), S => resultFA34, Cout => carryOutFA34);
FA35:full_adder port map (A => pp_ext(5)(30), B => pp_ext(6)(28), Cin => pp_ext(7)(26), S => resultFA35, Cout => carryOutFA35);
HA9:half_adder port map (A => pp_ext(8)(24), B => pp_ext(9)(22), S => resultHA9, Cout => carryOutHA9);
FA36:full_adder port map (A => pp_ext(3)(35), B => pp_ext(4)(33), Cin => pp_ext(5)(31), S => resultFA36, Cout => carryOutFA36);
FA37:full_adder port map (A => pp_ext(6)(29), B => pp_ext(7)(27), Cin => pp_ext(8)(25), S => resultFA37, Cout => carryOutFA37);
FA38:full_adder port map (A => pp_ext(3)(36), B => pp_ext(4)(34), Cin => pp_ext(5)(32), S => resultFA38, Cout => carryOutFA38);
HA10:half_adder port map (A => pp_ext(6)(30), B => pp_ext(7)(28), S => resultHA10, Cout => carryOutHA10);
FA39:full_adder port map (A => pp_ext(4)(35), B => pp_ext(5)(33), Cin => pp_ext(6)(31), S => resultFA39, Cout => carryOutFA39);
HA11:half_adder port map (A => pp_ext(4)(36), B => pp_ext(5)(34), S => resultHA11, Cout => carryOutHA11);
HA12:half_adder port map (A => pp_ext(0)(16), B => pp_ext(1)(16), S => resultHA12, Cout => carryOutHA12);
HA13:half_adder port map (A => pp_ext(0)(17), B => pp_ext(1)(17), S => resultHA13, Cout => carryOutHA13);
FA40:full_adder port map (A => pp_ext(0)(18), B => pp_ext(1)(18), Cin => pp_ext(2)(16), S => resultFA40, Cout => carryOutFA40);
HA14:half_adder port map (A => pp_ext(3)(14), B => pp_ext(4)(12), S => resultHA14, Cout => carryOutHA14);
FA41:full_adder port map (A => pp_ext(0)(19), B => pp_ext(1)(19), Cin => pp_ext(2)(17), S => resultFA41, Cout => carryOutFA41);
HA15:half_adder port map (A => pp_ext(3)(15), B => pp_ext(4)(13), S => resultHA15, Cout => carryOutHA15);
FA42:full_adder port map (A => pp_ext(0)(20), B => pp_ext(1)(20), Cin => pp_ext(2)(18), S => resultFA42, Cout => carryOutFA42);
FA43:full_adder port map (A => pp_ext(3)(16), B => pp_ext(4)(14), Cin => pp_ext(5)(12), S => resultFA43, Cout => carryOutFA43);
HA16:half_adder port map (A => pp_ext(6)(10), B => pp_ext(7)(8), S => resultHA16, Cout => carryOutHA16);
FA44:full_adder port map (A => pp_ext(0)(21), B => pp_ext(1)(21), Cin => pp_ext(2)(19), S => resultFA44, Cout => carryOutFA44);
FA45:full_adder port map (A => pp_ext(3)(17), B => pp_ext(4)(15), Cin => pp_ext(5)(13), S => resultFA45, Cout => carryOutFA45);
HA17:half_adder port map (A => pp_ext(6)(11), B => pp_ext(7)(9), S => resultHA17, Cout => carryOutHA17);
FA46:full_adder port map (A => pp_ext(0)(22), B => pp_ext(1)(22), Cin => pp_ext(2)(20), S => resultFA46, Cout => carryOutFA46);
FA47:full_adder port map (A => pp_ext(3)(18), B => pp_ext(4)(16), Cin => pp_ext(5)(14), S => resultFA47, Cout => carryOutFA47);
FA48:full_adder port map (A => pp_ext(6)(12), B => pp_ext(7)(10), Cin => pp_ext(8)(8), S => resultFA48, Cout => carryOutFA48);
HA18:half_adder port map (A => pp_ext(9)(6), B => pp_ext(10)(4), S => resultHA18, Cout => carryOutHA18);
FA49:full_adder port map (A => pp_ext(0)(23), B => pp_ext(1)(23), Cin => pp_ext(2)(21), S => resultFA49, Cout => carryOutFA49);
FA50:full_adder port map (A => pp_ext(3)(19), B => pp_ext(4)(17), Cin => pp_ext(5)(15), S => resultFA50, Cout => carryOutFA50);
FA51:full_adder port map (A => pp_ext(6)(13), B => pp_ext(7)(11), Cin => pp_ext(8)(9), S => resultFA51, Cout => carryOutFA51);
HA19:half_adder port map (A => pp_ext(9)(7), B => pp_ext(10)(5), S => resultHA19, Cout => carryOutHA19);
FA52:full_adder port map (A => resultHA0, B => pp_ext(2)(22), Cin => pp_ext(3)(20), S => resultFA52, Cout => carryOutFA52);
FA53:full_adder port map (A => pp_ext(4)(18), B => pp_ext(5)(16), Cin => pp_ext(6)(14), S => resultFA53, Cout => carryOutFA53);
FA54:full_adder port map (A => pp_ext(7)(12), B => pp_ext(8)(10), Cin => pp_ext(9)(8), S => resultFA54, Cout => carryOutFA54);
FA55:full_adder port map (A => pp_ext(10)(6), B => pp_ext(11)(4), Cin => pp_ext(12)(2), S => resultFA55, Cout => carryOutFA55);
FA56:full_adder port map (A => carryOutHA0, B => resultHA1, Cin => pp_ext(2)(23), S => resultFA56, Cout => carryOutFA56);
FA57:full_adder port map (A => pp_ext(3)(21), B => pp_ext(4)(19), Cin => pp_ext(5)(17), S => resultFA57, Cout => carryOutFA57);
FA58:full_adder port map (A => pp_ext(6)(15), B => pp_ext(7)(13), Cin => pp_ext(8)(11), S => resultFA58, Cout => carryOutFA58);
FA59:full_adder port map (A => pp_ext(9)(9), B => pp_ext(10)(7), Cin => pp_ext(11)(5), S => resultFA59, Cout => carryOutFA59);
FA60:full_adder port map (A => carryOutHA1, B => resultFA0, Cin => resultHA2, S => resultFA60, Cout => carryOutFA60);
FA61:full_adder port map (A => pp_ext(5)(18), B => pp_ext(6)(16), Cin => pp_ext(7)(14), S => resultFA61, Cout => carryOutFA61);
FA62:full_adder port map (A => pp_ext(8)(12), B => pp_ext(9)(10), Cin => pp_ext(10)(8), S => resultFA62, Cout => carryOutFA62);
FA63:full_adder port map (A => pp_ext(11)(6), B => pp_ext(12)(4), Cin => pp_ext(13)(2), S => resultFA63, Cout => carryOutFA63);
FA64:full_adder port map (A => carryOutFA0, B => carryOutHA2, Cin => resultFA1, S => resultFA64, Cout => carryOutFA64);
FA65:full_adder port map (A => resultHA3, B => pp_ext(5)(19), Cin => pp_ext(6)(17), S => resultFA65, Cout => carryOutFA65);
FA66:full_adder port map (A => pp_ext(7)(15), B => pp_ext(8)(13), Cin => pp_ext(9)(11), S => resultFA66, Cout => carryOutFA66);
FA67:full_adder port map (A => pp_ext(10)(9), B => pp_ext(11)(7), Cin => pp_ext(12)(5), S => resultFA67, Cout => carryOutFA67);
FA68:full_adder port map (A => carryOutFA1, B => carryOutHA3, Cin => resultFA2, S => resultFA68, Cout => carryOutFA68);
FA69:full_adder port map (A => resultFA3, B => resultHA4, Cin => pp_ext(8)(14), S => resultFA69, Cout => carryOutFA69);
FA70:full_adder port map (A => pp_ext(9)(12), B => pp_ext(10)(10), Cin => pp_ext(11)(8), S => resultFA70, Cout => carryOutFA70);
FA71:full_adder port map (A => pp_ext(12)(6), B => pp_ext(13)(4), Cin => pp_ext(14)(2), S => resultFA71, Cout => carryOutFA71);
FA72:full_adder port map (A => carryOutFA2, B => carryOutFA3, Cin => carryOutHA4, S => resultFA72, Cout => carryOutFA72);
FA73:full_adder port map (A => resultFA4, B => resultFA5, Cin => resultHA5, S => resultFA73, Cout => carryOutFA73);
FA74:full_adder port map (A => pp_ext(8)(15), B => pp_ext(9)(13), Cin => pp_ext(10)(11), S => resultFA74, Cout => carryOutFA74);
FA75:full_adder port map (A => pp_ext(11)(9), B => pp_ext(12)(7), Cin => pp_ext(13)(5), S => resultFA75, Cout => carryOutFA75);
FA76:full_adder port map (A => carryOutFA4, B => carryOutFA5, Cin => carryOutHA5, S => resultFA76, Cout => carryOutFA76);
FA77:full_adder port map (A => resultFA6, B => resultFA7, Cin => resultFA8, S => resultFA77, Cout => carryOutFA77);
FA78:full_adder port map (A => resultHA6, B => pp_ext(11)(10), Cin => pp_ext(12)(8), S => resultFA78, Cout => carryOutFA78);
FA79:full_adder port map (A => pp_ext(13)(6), B => pp_ext(14)(4), Cin => pp_ext(15)(2), S => resultFA79, Cout => carryOutFA79);
FA80:full_adder port map (A => carryOutFA6, B => carryOutFA7, Cin => carryOutFA8, S => resultFA80, Cout => carryOutFA80);
FA81:full_adder port map (A => carryOutHA6, B => resultFA9, Cin => resultFA10, S => resultFA81, Cout => carryOutFA81);
FA82:full_adder port map (A => resultFA11, B => resultHA7, Cin => pp_ext(11)(11), S => resultFA82, Cout => carryOutFA82);
FA83:full_adder port map (A => pp_ext(12)(9), B => pp_ext(13)(7), Cin => pp_ext(14)(5), S => resultFA83, Cout => carryOutFA83);
FA84:full_adder port map (A => carryOutFA9, B => carryOutFA10, Cin => carryOutFA11, S => resultFA84, Cout => carryOutFA84);
FA85:full_adder port map (A => carryOutHA7, B => resultFA12, Cin => resultFA13, S => resultFA85, Cout => carryOutFA85);
FA86:full_adder port map (A => resultFA14, B => resultFA15, Cin => pp_ext(12)(10), S => resultFA86, Cout => carryOutFA86);
FA87:full_adder port map (A => pp_ext(13)(8), B => pp_ext(14)(6), Cin => pp_ext(15)(4), S => resultFA87, Cout => carryOutFA87);
FA88:full_adder port map (A => carryOutFA12, B => carryOutFA13, Cin => carryOutFA14, S => resultFA88, Cout => carryOutFA88);
FA89:full_adder port map (A => carryOutFA15, B => resultFA16, Cin => resultFA17, S => resultFA89, Cout => carryOutFA89);
FA90:full_adder port map (A => resultFA18, B => resultFA19, Cin => pp_ext(12)(11), S => resultFA90, Cout => carryOutFA90);
FA91:full_adder port map (A => pp_ext(13)(9), B => pp_ext(14)(7), Cin => pp_ext(15)(5), S => resultFA91, Cout => carryOutFA91);
FA92:full_adder port map (A => carryOutFA16, B => carryOutFA17, Cin => carryOutFA18, S => resultFA92, Cout => carryOutFA92);
FA93:full_adder port map (A => carryOutFA19, B => resultFA20, Cin => resultFA21, S => resultFA93, Cout => carryOutFA93);
FA94:full_adder port map (A => resultFA22, B => resultFA23, Cin => pp_ext(12)(12), S => resultFA94, Cout => carryOutFA94);
FA95:full_adder port map (A => pp_ext(13)(10), B => pp_ext(14)(8), Cin => pp_ext(15)(6), S => resultFA95, Cout => carryOutFA95);
FA96:full_adder port map (A => carryOutFA20, B => carryOutFA21, Cin => carryOutFA22, S => resultFA96, Cout => carryOutFA96);
FA97:full_adder port map (A => carryOutFA23, B => resultFA24, Cin => resultFA25, S => resultFA97, Cout => carryOutFA97);
FA98:full_adder port map (A => resultFA26, B => resultFA27, Cin => pp_ext(12)(13), S => resultFA98, Cout => carryOutFA98);
FA99:full_adder port map (A => pp_ext(13)(11), B => pp_ext(14)(9), Cin => pp_ext(15)(7), S => resultFA99, Cout => carryOutFA99);
FA100:full_adder port map (A => carryOutFA24, B => carryOutFA25, Cin => carryOutFA26, S => resultFA100, Cout => carryOutFA100);
FA101:full_adder port map (A => carryOutFA27, B => resultFA28, Cin => resultFA29, S => resultFA101, Cout => carryOutFA101);
FA102:full_adder port map (A => resultFA30, B => resultHA8, Cin => pp_ext(12)(14), S => resultFA102, Cout => carryOutFA102);
FA103:full_adder port map (A => pp_ext(13)(12), B => pp_ext(14)(10), Cin => pp_ext(15)(8), S => resultFA103, Cout => carryOutFA103);
FA104:full_adder port map (A => carryOutFA28, B => carryOutFA29, Cin => carryOutFA30, S => resultFA104, Cout => carryOutFA104);
FA105:full_adder port map (A => carryOutHA8, B => resultFA31, Cin => resultFA32, S => resultFA105, Cout => carryOutFA105);
FA106:full_adder port map (A => resultFA33, B => pp_ext(11)(17), Cin => pp_ext(12)(15), S => resultFA106, Cout => carryOutFA106);
FA107:full_adder port map (A => pp_ext(13)(13), B => pp_ext(14)(11), Cin => pp_ext(15)(9), S => resultFA107, Cout => carryOutFA107);
FA108:full_adder port map (A => carryOutFA31, B => carryOutFA32, Cin => carryOutFA33, S => resultFA108, Cout => carryOutFA108);
FA109:full_adder port map (A => resultFA34, B => resultFA35, Cin => resultHA9, S => resultFA109, Cout => carryOutFA109);
FA110:full_adder port map (A => pp_ext(10)(20), B => pp_ext(11)(18), Cin => pp_ext(12)(16), S => resultFA110, Cout => carryOutFA110);
FA111:full_adder port map (A => pp_ext(13)(14), B => pp_ext(14)(12), Cin => pp_ext(15)(10), S => resultFA111, Cout => carryOutFA111);
FA112:full_adder port map (A => carryOutFA34, B => carryOutFA35, Cin => carryOutHA9, S => resultFA112, Cout => carryOutFA112);
FA113:full_adder port map (A => resultFA36, B => resultFA37, Cin => pp_ext(9)(23), S => resultFA113, Cout => carryOutFA113);
FA114:full_adder port map (A => pp_ext(10)(21), B => pp_ext(11)(19), Cin => pp_ext(12)(17), S => resultFA114, Cout => carryOutFA114);
FA115:full_adder port map (A => pp_ext(13)(15), B => pp_ext(14)(13), Cin => pp_ext(15)(11), S => resultFA115, Cout => carryOutFA115);
FA116:full_adder port map (A => carryOutFA36, B => carryOutFA37, Cin => resultFA38, S => resultFA116, Cout => carryOutFA116);
FA117:full_adder port map (A => resultHA10, B => pp_ext(8)(26), Cin => pp_ext(9)(24), S => resultFA117, Cout => carryOutFA117);
FA118:full_adder port map (A => pp_ext(10)(22), B => pp_ext(11)(20), Cin => pp_ext(12)(18), S => resultFA118, Cout => carryOutFA118);
FA119:full_adder port map (A => pp_ext(13)(16), B => pp_ext(14)(14), Cin => pp_ext(15)(12), S => resultFA119, Cout => carryOutFA119);
FA120:full_adder port map (A => carryOutFA38, B => carryOutHA10, Cin => resultFA39, S => resultFA120, Cout => carryOutFA120);
FA121:full_adder port map (A => pp_ext(7)(29), B => pp_ext(8)(27), Cin => pp_ext(9)(25), S => resultFA121, Cout => carryOutFA121);
FA122:full_adder port map (A => pp_ext(10)(23), B => pp_ext(11)(21), Cin => pp_ext(12)(19), S => resultFA122, Cout => carryOutFA122);
FA123:full_adder port map (A => pp_ext(13)(17), B => pp_ext(14)(15), Cin => pp_ext(15)(13), S => resultFA123, Cout => carryOutFA123);
FA124:full_adder port map (A => carryOutFA39, B => resultHA11, Cin => pp_ext(6)(32), S => resultFA124, Cout => carryOutFA124);
FA125:full_adder port map (A => pp_ext(7)(30), B => pp_ext(8)(28), Cin => pp_ext(9)(26), S => resultFA125, Cout => carryOutFA125);
FA126:full_adder port map (A => pp_ext(10)(24), B => pp_ext(11)(22), Cin => pp_ext(12)(20), S => resultFA126, Cout => carryOutFA126);
FA127:full_adder port map (A => pp_ext(13)(18), B => pp_ext(14)(16), Cin => pp_ext(15)(14), S => resultFA127, Cout => carryOutFA127);
FA128:full_adder port map (A => carryOutHA11, B => pp_ext(5)(35), Cin => pp_ext(6)(33), S => resultFA128, Cout => carryOutFA128);
FA129:full_adder port map (A => pp_ext(7)(31), B => pp_ext(8)(29), Cin => pp_ext(9)(27), S => resultFA129, Cout => carryOutFA129);
FA130:full_adder port map (A => pp_ext(10)(25), B => pp_ext(11)(23), Cin => pp_ext(12)(21), S => resultFA130, Cout => carryOutFA130);
FA131:full_adder port map (A => pp_ext(13)(19), B => pp_ext(14)(17), Cin => pp_ext(15)(15), S => resultFA131, Cout => carryOutFA131);
FA132:full_adder port map (A => pp_ext(5)(36), B => pp_ext(6)(34), Cin => pp_ext(7)(32), S => resultFA132, Cout => carryOutFA132);
FA133:full_adder port map (A => pp_ext(8)(30), B => pp_ext(9)(28), Cin => pp_ext(10)(26), S => resultFA133, Cout => carryOutFA133);
FA134:full_adder port map (A => pp_ext(11)(24), B => pp_ext(12)(22), Cin => pp_ext(13)(20), S => resultFA134, Cout => carryOutFA134);
HA20:half_adder port map (A => pp_ext(14)(18), B => pp_ext(15)(16), S => resultHA20, Cout => carryOutHA20);
FA135:full_adder port map (A => pp_ext(6)(35), B => pp_ext(7)(33), Cin => pp_ext(8)(31), S => resultFA135, Cout => carryOutFA135);
FA136:full_adder port map (A => pp_ext(9)(29), B => pp_ext(10)(27), Cin => pp_ext(11)(25), S => resultFA136, Cout => carryOutFA136);
FA137:full_adder port map (A => pp_ext(12)(23), B => pp_ext(13)(21), Cin => pp_ext(14)(19), S => resultFA137, Cout => carryOutFA137);
FA138:full_adder port map (A => pp_ext(6)(36), B => pp_ext(7)(34), Cin => pp_ext(8)(32), S => resultFA138, Cout => carryOutFA138);
FA139:full_adder port map (A => pp_ext(9)(30), B => pp_ext(10)(28), Cin => pp_ext(11)(26), S => resultFA139, Cout => carryOutFA139);
HA21:half_adder port map (A => pp_ext(12)(24), B => pp_ext(13)(22), S => resultHA21, Cout => carryOutHA21);
FA140:full_adder port map (A => pp_ext(7)(35), B => pp_ext(8)(33), Cin => pp_ext(9)(31), S => resultFA140, Cout => carryOutFA140);
FA141:full_adder port map (A => pp_ext(10)(29), B => pp_ext(11)(27), Cin => pp_ext(12)(25), S => resultFA141, Cout => carryOutFA141);
FA142:full_adder port map (A => pp_ext(7)(36), B => pp_ext(8)(34), Cin => pp_ext(9)(32), S => resultFA142, Cout => carryOutFA142);
HA22:half_adder port map (A => pp_ext(10)(30), B => pp_ext(11)(28), S => resultHA22, Cout => carryOutHA22);
FA143:full_adder port map (A => pp_ext(8)(35), B => pp_ext(9)(33), Cin => pp_ext(10)(31), S => resultFA143, Cout => carryOutFA143);
HA23:half_adder port map (A => pp_ext(8)(36), B => pp_ext(9)(34), S => resultHA23, Cout => carryOutHA23);
HA24:half_adder port map (A => pp_ext(0)(10), B => pp_ext(1)(10), S => resultHA24, Cout => carryOutHA24);
HA25:half_adder port map (A => pp_ext(0)(11), B => pp_ext(1)(11), S => resultHA25, Cout => carryOutHA25);
FA144:full_adder port map (A => pp_ext(0)(12), B => pp_ext(1)(12), Cin => pp_ext(2)(10), S => resultFA144, Cout => carryOutFA144);
HA26:half_adder port map (A => pp_ext(3)(8), B => pp_ext(4)(6), S => resultHA26, Cout => carryOutHA26);
FA145:full_adder port map (A => pp_ext(0)(13), B => pp_ext(1)(13), Cin => pp_ext(2)(11), S => resultFA145, Cout => carryOutFA145);
HA27:half_adder port map (A => pp_ext(3)(9), B => pp_ext(4)(7), S => resultHA27, Cout => carryOutHA27);
FA146:full_adder port map (A => pp_ext(0)(14), B => pp_ext(1)(14), Cin => pp_ext(2)(12), S => resultFA146, Cout => carryOutFA146);
FA147:full_adder port map (A => pp_ext(3)(10), B => pp_ext(4)(8), Cin => pp_ext(5)(6), S => resultFA147, Cout => carryOutFA147);
HA28:half_adder port map (A => pp_ext(6)(4), B => pp_ext(7)(2), S => resultHA28, Cout => carryOutHA28);
FA148:full_adder port map (A => pp_ext(0)(15), B => pp_ext(1)(15), Cin => pp_ext(2)(13), S => resultFA148, Cout => carryOutFA148);
FA149:full_adder port map (A => pp_ext(3)(11), B => pp_ext(4)(9), Cin => pp_ext(5)(7), S => resultFA149, Cout => carryOutFA149);
HA29:half_adder port map (A => pp_ext(6)(5), B => pp_ext(7)(3), S => resultHA29, Cout => carryOutHA29);
FA150:full_adder port map (A => resultHA12, B => pp_ext(2)(14), Cin => pp_ext(3)(12), S => resultFA150, Cout => carryOutFA150);
FA151:full_adder port map (A => pp_ext(4)(10), B => pp_ext(5)(8), Cin => pp_ext(6)(6), S => resultFA151, Cout => carryOutFA151);
FA152:full_adder port map (A => pp_ext(7)(4), B => pp_ext(8)(2), Cin => pp_ext(9)(0), S => resultFA152, Cout => carryOutFA152);
FA153:full_adder port map (A => carryOutHA12, B => resultHA13, Cin => pp_ext(2)(15), S => resultFA153, Cout => carryOutFA153);
FA154:full_adder port map (A => pp_ext(3)(13), B => pp_ext(4)(11), Cin => pp_ext(5)(9), S => resultFA154, Cout => carryOutFA154);
FA155:full_adder port map (A => pp_ext(6)(7), B => pp_ext(7)(5), Cin => pp_ext(8)(3), S => resultFA155, Cout => carryOutFA155);
FA156:full_adder port map (A => carryOutHA13, B => resultFA40, Cin => resultHA14, S => resultFA156, Cout => carryOutFA156);
FA157:full_adder port map (A => pp_ext(5)(10), B => pp_ext(6)(8), Cin => pp_ext(7)(6), S => resultFA157, Cout => carryOutFA157);
FA158:full_adder port map (A => pp_ext(8)(4), B => pp_ext(9)(2), Cin => pp_ext(10)(0), S => resultFA158, Cout => carryOutFA158);
FA159:full_adder port map (A => carryOutFA40, B => carryOutHA14, Cin => resultFA41, S => resultFA159, Cout => carryOutFA159);
FA160:full_adder port map (A => resultHA15, B => pp_ext(5)(11), Cin => pp_ext(6)(9), S => resultFA160, Cout => carryOutFA160);
FA161:full_adder port map (A => pp_ext(7)(7), B => pp_ext(8)(5), Cin => pp_ext(9)(3), S => resultFA161, Cout => carryOutFA161);
FA162:full_adder port map (A => carryOutFA41, B => carryOutHA15, Cin => resultFA42, S => resultFA162, Cout => carryOutFA162);
FA163:full_adder port map (A => resultFA43, B => resultHA16, Cin => pp_ext(8)(6), S => resultFA163, Cout => carryOutFA163);
FA164:full_adder port map (A => pp_ext(9)(4), B => pp_ext(10)(2), Cin => pp_ext(11)(0), S => resultFA164, Cout => carryOutFA164);
FA165:full_adder port map (A => carryOutFA42, B => carryOutFA43, Cin => carryOutHA16, S => resultFA165, Cout => carryOutFA165);
FA166:full_adder port map (A => resultFA44, B => resultFA45, Cin => resultHA17, S => resultFA166, Cout => carryOutFA166);
FA167:full_adder port map (A => pp_ext(8)(7), B => pp_ext(9)(5), Cin => pp_ext(10)(3), S => resultFA167, Cout => carryOutFA167);
FA168:full_adder port map (A => carryOutFA44, B => carryOutFA45, Cin => carryOutHA17, S => resultFA168, Cout => carryOutFA168);
FA169:full_adder port map (A => resultFA46, B => resultFA47, Cin => resultFA48, S => resultFA169, Cout => carryOutFA169);
FA170:full_adder port map (A => resultHA18, B => pp_ext(11)(2), Cin => pp_ext(12)(0), S => resultFA170, Cout => carryOutFA170);
FA171:full_adder port map (A => carryOutFA46, B => carryOutFA47, Cin => carryOutFA48, S => resultFA171, Cout => carryOutFA171);
FA172:full_adder port map (A => carryOutHA18, B => resultFA49, Cin => resultFA50, S => resultFA172, Cout => carryOutFA172);
FA173:full_adder port map (A => resultFA51, B => resultHA19, Cin => pp_ext(11)(3), S => resultFA173, Cout => carryOutFA173);
FA174:full_adder port map (A => carryOutFA49, B => carryOutFA50, Cin => carryOutFA51, S => resultFA174, Cout => carryOutFA174);
FA175:full_adder port map (A => carryOutHA19, B => resultFA52, Cin => resultFA53, S => resultFA175, Cout => carryOutFA175);
FA176:full_adder port map (A => resultFA54, B => resultFA55, Cin => pp_ext(13)(0), S => resultFA176, Cout => carryOutFA176);
FA177:full_adder port map (A => carryOutFA52, B => carryOutFA53, Cin => carryOutFA54, S => resultFA177, Cout => carryOutFA177);
FA178:full_adder port map (A => carryOutFA55, B => resultFA56, Cin => resultFA57, S => resultFA178, Cout => carryOutFA178);
FA179:full_adder port map (A => resultFA58, B => resultFA59, Cin => pp_ext(12)(3), S => resultFA179, Cout => carryOutFA179);
FA180:full_adder port map (A => carryOutFA56, B => carryOutFA57, Cin => carryOutFA58, S => resultFA180, Cout => carryOutFA180);
FA181:full_adder port map (A => carryOutFA59, B => resultFA60, Cin => resultFA61, S => resultFA181, Cout => carryOutFA181);
FA182:full_adder port map (A => resultFA62, B => resultFA63, Cin => pp_ext(14)(0), S => resultFA182, Cout => carryOutFA182);
FA183:full_adder port map (A => carryOutFA60, B => carryOutFA61, Cin => carryOutFA62, S => resultFA183, Cout => carryOutFA183);
FA184:full_adder port map (A => carryOutFA63, B => resultFA64, Cin => resultFA65, S => resultFA184, Cout => carryOutFA184);
FA185:full_adder port map (A => resultFA66, B => resultFA67, Cin => pp_ext(13)(3), S => resultFA185, Cout => carryOutFA185);
FA186:full_adder port map (A => carryOutFA64, B => carryOutFA65, Cin => carryOutFA66, S => resultFA186, Cout => carryOutFA186);
FA187:full_adder port map (A => carryOutFA67, B => resultFA68, Cin => resultFA69, S => resultFA187, Cout => carryOutFA187);
FA188:full_adder port map (A => resultFA70, B => resultFA71, Cin => pp_ext(15)(0), S => resultFA188, Cout => carryOutFA188);
FA189:full_adder port map (A => carryOutFA68, B => carryOutFA69, Cin => carryOutFA70, S => resultFA189, Cout => carryOutFA189);
FA190:full_adder port map (A => carryOutFA71, B => resultFA72, Cin => resultFA73, S => resultFA190, Cout => carryOutFA190);
FA191:full_adder port map (A => resultFA74, B => resultFA75, Cin => pp_ext(14)(3), S => resultFA191, Cout => carryOutFA191);
FA192:full_adder port map (A => carryOutFA72, B => carryOutFA73, Cin => carryOutFA74, S => resultFA192, Cout => carryOutFA192);
FA193:full_adder port map (A => carryOutFA75, B => resultFA76, Cin => resultFA77, S => resultFA193, Cout => carryOutFA193);
FA194:full_adder port map (A => resultFA78, B => resultFA79, Cin => pp_ext(16)(0), S => resultFA194, Cout => carryOutFA194);
FA195:full_adder port map (A => carryOutFA76, B => carryOutFA77, Cin => carryOutFA78, S => resultFA195, Cout => carryOutFA195);
FA196:full_adder port map (A => carryOutFA79, B => resultFA80, Cin => resultFA81, S => resultFA196, Cout => carryOutFA196);
FA197:full_adder port map (A => resultFA82, B => resultFA83, Cin => pp_ext(15)(3), S => resultFA197, Cout => carryOutFA197);
FA198:full_adder port map (A => carryOutFA80, B => carryOutFA81, Cin => carryOutFA82, S => resultFA198, Cout => carryOutFA198);
FA199:full_adder port map (A => carryOutFA83, B => resultFA84, Cin => resultFA85, S => resultFA199, Cout => carryOutFA199);
FA200:full_adder port map (A => resultFA86, B => resultFA87, Cin => pp_ext(16)(2), S => resultFA200, Cout => carryOutFA200);
FA201:full_adder port map (A => carryOutFA84, B => carryOutFA85, Cin => carryOutFA86, S => resultFA201, Cout => carryOutFA201);
FA202:full_adder port map (A => carryOutFA87, B => resultFA88, Cin => resultFA89, S => resultFA202, Cout => carryOutFA202);
FA203:full_adder port map (A => resultFA90, B => resultFA91, Cin => pp_ext(16)(3), S => resultFA203, Cout => carryOutFA203);
FA204:full_adder port map (A => carryOutFA88, B => carryOutFA89, Cin => carryOutFA90, S => resultFA204, Cout => carryOutFA204);
FA205:full_adder port map (A => carryOutFA91, B => resultFA92, Cin => resultFA93, S => resultFA205, Cout => carryOutFA205);
FA206:full_adder port map (A => resultFA94, B => resultFA95, Cin => pp_ext(16)(4), S => resultFA206, Cout => carryOutFA206);
FA207:full_adder port map (A => carryOutFA92, B => carryOutFA93, Cin => carryOutFA94, S => resultFA207, Cout => carryOutFA207);
FA208:full_adder port map (A => carryOutFA95, B => resultFA96, Cin => resultFA97, S => resultFA208, Cout => carryOutFA208);
FA209:full_adder port map (A => resultFA98, B => resultFA99, Cin => pp_ext(16)(5), S => resultFA209, Cout => carryOutFA209);
FA210:full_adder port map (A => carryOutFA96, B => carryOutFA97, Cin => carryOutFA98, S => resultFA210, Cout => carryOutFA210);
FA211:full_adder port map (A => carryOutFA99, B => resultFA100, Cin => resultFA101, S => resultFA211, Cout => carryOutFA211);
FA212:full_adder port map (A => resultFA102, B => resultFA103, Cin => pp_ext(16)(6), S => resultFA212, Cout => carryOutFA212);
FA213:full_adder port map (A => carryOutFA100, B => carryOutFA101, Cin => carryOutFA102, S => resultFA213, Cout => carryOutFA213);
FA214:full_adder port map (A => carryOutFA103, B => resultFA104, Cin => resultFA105, S => resultFA214, Cout => carryOutFA214);
FA215:full_adder port map (A => resultFA106, B => resultFA107, Cin => pp_ext(16)(7), S => resultFA215, Cout => carryOutFA215);
FA216:full_adder port map (A => carryOutFA104, B => carryOutFA105, Cin => carryOutFA106, S => resultFA216, Cout => carryOutFA216);
FA217:full_adder port map (A => carryOutFA107, B => resultFA108, Cin => resultFA109, S => resultFA217, Cout => carryOutFA217);
FA218:full_adder port map (A => resultFA110, B => resultFA111, Cin => pp_ext(16)(8), S => resultFA218, Cout => carryOutFA218);
FA219:full_adder port map (A => carryOutFA108, B => carryOutFA109, Cin => carryOutFA110, S => resultFA219, Cout => carryOutFA219);
FA220:full_adder port map (A => carryOutFA111, B => resultFA112, Cin => resultFA113, S => resultFA220, Cout => carryOutFA220);
FA221:full_adder port map (A => resultFA114, B => resultFA115, Cin => pp_ext(16)(9), S => resultFA221, Cout => carryOutFA221);
FA222:full_adder port map (A => carryOutFA112, B => carryOutFA113, Cin => carryOutFA114, S => resultFA222, Cout => carryOutFA222);
FA223:full_adder port map (A => carryOutFA115, B => resultFA116, Cin => resultFA117, S => resultFA223, Cout => carryOutFA223);
FA224:full_adder port map (A => resultFA118, B => resultFA119, Cin => pp_ext(16)(10), S => resultFA224, Cout => carryOutFA224);
FA225:full_adder port map (A => carryOutFA116, B => carryOutFA117, Cin => carryOutFA118, S => resultFA225, Cout => carryOutFA225);
FA226:full_adder port map (A => carryOutFA119, B => resultFA120, Cin => resultFA121, S => resultFA226, Cout => carryOutFA226);
FA227:full_adder port map (A => resultFA122, B => resultFA123, Cin => pp_ext(16)(11), S => resultFA227, Cout => carryOutFA227);
FA228:full_adder port map (A => carryOutFA120, B => carryOutFA121, Cin => carryOutFA122, S => resultFA228, Cout => carryOutFA228);
FA229:full_adder port map (A => carryOutFA123, B => resultFA124, Cin => resultFA125, S => resultFA229, Cout => carryOutFA229);
FA230:full_adder port map (A => resultFA126, B => resultFA127, Cin => pp_ext(16)(12), S => resultFA230, Cout => carryOutFA230);
FA231:full_adder port map (A => carryOutFA124, B => carryOutFA125, Cin => carryOutFA126, S => resultFA231, Cout => carryOutFA231);
FA232:full_adder port map (A => carryOutFA127, B => resultFA128, Cin => resultFA129, S => resultFA232, Cout => carryOutFA232);
FA233:full_adder port map (A => resultFA130, B => resultFA131, Cin => pp_ext(16)(13), S => resultFA233, Cout => carryOutFA233);
FA234:full_adder port map (A => carryOutFA128, B => carryOutFA129, Cin => carryOutFA130, S => resultFA234, Cout => carryOutFA234);
FA235:full_adder port map (A => carryOutFA131, B => resultFA132, Cin => resultFA133, S => resultFA235, Cout => carryOutFA235);
FA236:full_adder port map (A => resultFA134, B => resultHA20, Cin => pp_ext(16)(14), S => resultFA236, Cout => carryOutFA236);
FA237:full_adder port map (A => carryOutFA132, B => carryOutFA133, Cin => carryOutFA134, S => resultFA237, Cout => carryOutFA237);
FA238:full_adder port map (A => carryOutHA20, B => resultFA135, Cin => resultFA136, S => resultFA238, Cout => carryOutFA238);
FA239:full_adder port map (A => resultFA137, B => pp_ext(15)(17), Cin => pp_ext(16)(15), S => resultFA239, Cout => carryOutFA239);
FA240:full_adder port map (A => carryOutFA135, B => carryOutFA136, Cin => carryOutFA137, S => resultFA240, Cout => carryOutFA240);
FA241:full_adder port map (A => resultFA138, B => resultFA139, Cin => resultHA21, S => resultFA241, Cout => carryOutFA241);
FA242:full_adder port map (A => pp_ext(14)(20), B => pp_ext(15)(18), Cin => pp_ext(16)(16), S => resultFA242, Cout => carryOutFA242);
FA243:full_adder port map (A => carryOutFA138, B => carryOutFA139, Cin => carryOutHA21, S => resultFA243, Cout => carryOutFA243);
FA244:full_adder port map (A => resultFA140, B => resultFA141, Cin => pp_ext(13)(23), S => resultFA244, Cout => carryOutFA244);
FA245:full_adder port map (A => pp_ext(14)(21), B => pp_ext(15)(19), Cin => pp_ext(16)(17), S => resultFA245, Cout => carryOutFA245);
FA246:full_adder port map (A => carryOutFA140, B => carryOutFA141, Cin => resultFA142, S => resultFA246, Cout => carryOutFA246);
FA247:full_adder port map (A => resultHA22, B => pp_ext(12)(26), Cin => pp_ext(13)(24), S => resultFA247, Cout => carryOutFA247);
FA248:full_adder port map (A => pp_ext(14)(22), B => pp_ext(15)(20), Cin => pp_ext(16)(18), S => resultFA248, Cout => carryOutFA248);
FA249:full_adder port map (A => carryOutFA142, B => carryOutHA22, Cin => resultFA143, S => resultFA249, Cout => carryOutFA249);
FA250:full_adder port map (A => pp_ext(11)(29), B => pp_ext(12)(27), Cin => pp_ext(13)(25), S => resultFA250, Cout => carryOutFA250);
FA251:full_adder port map (A => pp_ext(14)(23), B => pp_ext(15)(21), Cin => pp_ext(16)(19), S => resultFA251, Cout => carryOutFA251);
FA252:full_adder port map (A => carryOutFA143, B => resultHA23, Cin => pp_ext(10)(32), S => resultFA252, Cout => carryOutFA252);
FA253:full_adder port map (A => pp_ext(11)(30), B => pp_ext(12)(28), Cin => pp_ext(13)(26), S => resultFA253, Cout => carryOutFA253);
FA254:full_adder port map (A => pp_ext(14)(24), B => pp_ext(15)(22), Cin => pp_ext(16)(20), S => resultFA254, Cout => carryOutFA254);
FA255:full_adder port map (A => carryOutHA23, B => pp_ext(9)(35), Cin => pp_ext(10)(33), S => resultFA255, Cout => carryOutFA255);
FA256:full_adder port map (A => pp_ext(11)(31), B => pp_ext(12)(29), Cin => pp_ext(13)(27), S => resultFA256, Cout => carryOutFA256);
FA257:full_adder port map (A => pp_ext(14)(25), B => pp_ext(15)(23), Cin => pp_ext(16)(21), S => resultFA257, Cout => carryOutFA257);
FA258:full_adder port map (A => pp_ext(9)(36), B => pp_ext(10)(34), Cin => pp_ext(11)(32), S => resultFA258, Cout => carryOutFA258);
FA259:full_adder port map (A => pp_ext(12)(30), B => pp_ext(13)(28), Cin => pp_ext(14)(26), S => resultFA259, Cout => carryOutFA259);
HA30:half_adder port map (A => pp_ext(15)(24), B => pp_ext(16)(22), S => resultHA30, Cout => carryOutHA30);
FA260:full_adder port map (A => pp_ext(10)(35), B => pp_ext(11)(33), Cin => pp_ext(12)(31), S => resultFA260, Cout => carryOutFA260);
FA261:full_adder port map (A => pp_ext(13)(29), B => pp_ext(14)(27), Cin => pp_ext(15)(25), S => resultFA261, Cout => carryOutFA261);
FA262:full_adder port map (A => pp_ext(10)(36), B => pp_ext(11)(34), Cin => pp_ext(12)(32), S => resultFA262, Cout => carryOutFA262);
HA31:half_adder port map (A => pp_ext(13)(30), B => pp_ext(14)(28), S => resultHA31, Cout => carryOutHA31);
FA263:full_adder port map (A => pp_ext(11)(35), B => pp_ext(12)(33), Cin => pp_ext(13)(31), S => resultFA263, Cout => carryOutFA263);
HA32:half_adder port map (A => pp_ext(11)(36), B => pp_ext(12)(34), S => resultHA32, Cout => carryOutHA32);
HA33:half_adder port map (A => pp_ext(0)(6), B => pp_ext(1)(6), S => resultHA33, Cout => carryOutHA33);
HA34:half_adder port map (A => pp_ext(0)(7), B => pp_ext(1)(7), S => resultHA34, Cout => carryOutHA34);
FA264:full_adder port map (A => pp_ext(0)(8), B => pp_ext(1)(8), Cin => pp_ext(2)(6), S => resultFA264, Cout => carryOutFA264);
HA35:half_adder port map (A => pp_ext(3)(4), B => pp_ext(4)(2), S => resultHA35, Cout => carryOutHA35);
FA265:full_adder port map (A => pp_ext(0)(9), B => pp_ext(1)(9), Cin => pp_ext(2)(7), S => resultFA265, Cout => carryOutFA265);
HA36:half_adder port map (A => pp_ext(3)(5), B => pp_ext(4)(3), S => resultHA36, Cout => carryOutHA36);
FA266:full_adder port map (A => resultHA24, B => pp_ext(2)(8), Cin => pp_ext(3)(6), S => resultFA266, Cout => carryOutFA266);
FA267:full_adder port map (A => pp_ext(4)(4), B => pp_ext(5)(2), Cin => pp_ext(6)(0), S => resultFA267, Cout => carryOutFA267);
FA268:full_adder port map (A => carryOutHA24, B => resultHA25, Cin => pp_ext(2)(9), S => resultFA268, Cout => carryOutFA268);
FA269:full_adder port map (A => pp_ext(3)(7), B => pp_ext(4)(5), Cin => pp_ext(5)(3), S => resultFA269, Cout => carryOutFA269);
FA270:full_adder port map (A => carryOutHA25, B => resultFA144, Cin => resultHA26, S => resultFA270, Cout => carryOutFA270);
FA271:full_adder port map (A => pp_ext(5)(4), B => pp_ext(6)(2), Cin => pp_ext(7)(0), S => resultFA271, Cout => carryOutFA271);
FA272:full_adder port map (A => carryOutFA144, B => carryOutHA26, Cin => resultFA145, S => resultFA272, Cout => carryOutFA272);
FA273:full_adder port map (A => resultHA27, B => pp_ext(5)(5), Cin => pp_ext(6)(3), S => resultFA273, Cout => carryOutFA273);
FA274:full_adder port map (A => carryOutFA145, B => carryOutHA27, Cin => resultFA146, S => resultFA274, Cout => carryOutFA274);
FA275:full_adder port map (A => resultFA147, B => resultHA28, Cin => pp_ext(8)(0), S => resultFA275, Cout => carryOutFA275);
FA276:full_adder port map (A => carryOutFA146, B => carryOutFA147, Cin => carryOutHA28, S => resultFA276, Cout => carryOutFA276);
FA277:full_adder port map (A => resultFA148, B => resultFA149, Cin => resultHA29, S => resultFA277, Cout => carryOutFA277);
FA278:full_adder port map (A => carryOutFA148, B => carryOutFA149, Cin => carryOutHA29, S => resultFA278, Cout => carryOutFA278);
FA279:full_adder port map (A => resultFA150, B => resultFA151, Cin => resultFA152, S => resultFA279, Cout => carryOutFA279);
FA280:full_adder port map (A => carryOutFA150, B => carryOutFA151, Cin => carryOutFA152, S => resultFA280, Cout => carryOutFA280);
FA281:full_adder port map (A => resultFA153, B => resultFA154, Cin => resultFA155, S => resultFA281, Cout => carryOutFA281);
FA282:full_adder port map (A => carryOutFA153, B => carryOutFA154, Cin => carryOutFA155, S => resultFA282, Cout => carryOutFA282);
FA283:full_adder port map (A => resultFA156, B => resultFA157, Cin => resultFA158, S => resultFA283, Cout => carryOutFA283);
FA284:full_adder port map (A => carryOutFA156, B => carryOutFA157, Cin => carryOutFA158, S => resultFA284, Cout => carryOutFA284);
FA285:full_adder port map (A => resultFA159, B => resultFA160, Cin => resultFA161, S => resultFA285, Cout => carryOutFA285);
FA286:full_adder port map (A => carryOutFA159, B => carryOutFA160, Cin => carryOutFA161, S => resultFA286, Cout => carryOutFA286);
FA287:full_adder port map (A => resultFA162, B => resultFA163, Cin => resultFA164, S => resultFA287, Cout => carryOutFA287);
FA288:full_adder port map (A => carryOutFA162, B => carryOutFA163, Cin => carryOutFA164, S => resultFA288, Cout => carryOutFA288);
FA289:full_adder port map (A => resultFA165, B => resultFA166, Cin => resultFA167, S => resultFA289, Cout => carryOutFA289);
FA290:full_adder port map (A => carryOutFA165, B => carryOutFA166, Cin => carryOutFA167, S => resultFA290, Cout => carryOutFA290);
FA291:full_adder port map (A => resultFA168, B => resultFA169, Cin => resultFA170, S => resultFA291, Cout => carryOutFA291);
FA292:full_adder port map (A => carryOutFA168, B => carryOutFA169, Cin => carryOutFA170, S => resultFA292, Cout => carryOutFA292);
FA293:full_adder port map (A => resultFA171, B => resultFA172, Cin => resultFA173, S => resultFA293, Cout => carryOutFA293);
FA294:full_adder port map (A => carryOutFA171, B => carryOutFA172, Cin => carryOutFA173, S => resultFA294, Cout => carryOutFA294);
FA295:full_adder port map (A => resultFA174, B => resultFA175, Cin => resultFA176, S => resultFA295, Cout => carryOutFA295);
FA296:full_adder port map (A => carryOutFA174, B => carryOutFA175, Cin => carryOutFA176, S => resultFA296, Cout => carryOutFA296);
FA297:full_adder port map (A => resultFA177, B => resultFA178, Cin => resultFA179, S => resultFA297, Cout => carryOutFA297);
FA298:full_adder port map (A => carryOutFA177, B => carryOutFA178, Cin => carryOutFA179, S => resultFA298, Cout => carryOutFA298);
FA299:full_adder port map (A => resultFA180, B => resultFA181, Cin => resultFA182, S => resultFA299, Cout => carryOutFA299);
FA300:full_adder port map (A => carryOutFA180, B => carryOutFA181, Cin => carryOutFA182, S => resultFA300, Cout => carryOutFA300);
FA301:full_adder port map (A => resultFA183, B => resultFA184, Cin => resultFA185, S => resultFA301, Cout => carryOutFA301);
FA302:full_adder port map (A => carryOutFA183, B => carryOutFA184, Cin => carryOutFA185, S => resultFA302, Cout => carryOutFA302);
FA303:full_adder port map (A => resultFA186, B => resultFA187, Cin => resultFA188, S => resultFA303, Cout => carryOutFA303);
FA304:full_adder port map (A => carryOutFA186, B => carryOutFA187, Cin => carryOutFA188, S => resultFA304, Cout => carryOutFA304);
FA305:full_adder port map (A => resultFA189, B => resultFA190, Cin => resultFA191, S => resultFA305, Cout => carryOutFA305);
FA306:full_adder port map (A => carryOutFA189, B => carryOutFA190, Cin => carryOutFA191, S => resultFA306, Cout => carryOutFA306);
FA307:full_adder port map (A => resultFA192, B => resultFA193, Cin => resultFA194, S => resultFA307, Cout => carryOutFA307);
FA308:full_adder port map (A => carryOutFA192, B => carryOutFA193, Cin => carryOutFA194, S => resultFA308, Cout => carryOutFA308);
FA309:full_adder port map (A => resultFA195, B => resultFA196, Cin => resultFA197, S => resultFA309, Cout => carryOutFA309);
FA310:full_adder port map (A => carryOutFA195, B => carryOutFA196, Cin => carryOutFA197, S => resultFA310, Cout => carryOutFA310);
FA311:full_adder port map (A => resultFA198, B => resultFA199, Cin => resultFA200, S => resultFA311, Cout => carryOutFA311);
FA312:full_adder port map (A => carryOutFA198, B => carryOutFA199, Cin => carryOutFA200, S => resultFA312, Cout => carryOutFA312);
FA313:full_adder port map (A => resultFA201, B => resultFA202, Cin => resultFA203, S => resultFA313, Cout => carryOutFA313);
FA314:full_adder port map (A => carryOutFA201, B => carryOutFA202, Cin => carryOutFA203, S => resultFA314, Cout => carryOutFA314);
FA315:full_adder port map (A => resultFA204, B => resultFA205, Cin => resultFA206, S => resultFA315, Cout => carryOutFA315);
FA316:full_adder port map (A => carryOutFA204, B => carryOutFA205, Cin => carryOutFA206, S => resultFA316, Cout => carryOutFA316);
FA317:full_adder port map (A => resultFA207, B => resultFA208, Cin => resultFA209, S => resultFA317, Cout => carryOutFA317);
FA318:full_adder port map (A => carryOutFA207, B => carryOutFA208, Cin => carryOutFA209, S => resultFA318, Cout => carryOutFA318);
FA319:full_adder port map (A => resultFA210, B => resultFA211, Cin => resultFA212, S => resultFA319, Cout => carryOutFA319);
FA320:full_adder port map (A => carryOutFA210, B => carryOutFA211, Cin => carryOutFA212, S => resultFA320, Cout => carryOutFA320);
FA321:full_adder port map (A => resultFA213, B => resultFA214, Cin => resultFA215, S => resultFA321, Cout => carryOutFA321);
FA322:full_adder port map (A => carryOutFA213, B => carryOutFA214, Cin => carryOutFA215, S => resultFA322, Cout => carryOutFA322);
FA323:full_adder port map (A => resultFA216, B => resultFA217, Cin => resultFA218, S => resultFA323, Cout => carryOutFA323);
FA324:full_adder port map (A => carryOutFA216, B => carryOutFA217, Cin => carryOutFA218, S => resultFA324, Cout => carryOutFA324);
FA325:full_adder port map (A => resultFA219, B => resultFA220, Cin => resultFA221, S => resultFA325, Cout => carryOutFA325);
FA326:full_adder port map (A => carryOutFA219, B => carryOutFA220, Cin => carryOutFA221, S => resultFA326, Cout => carryOutFA326);
FA327:full_adder port map (A => resultFA222, B => resultFA223, Cin => resultFA224, S => resultFA327, Cout => carryOutFA327);
FA328:full_adder port map (A => carryOutFA222, B => carryOutFA223, Cin => carryOutFA224, S => resultFA328, Cout => carryOutFA328);
FA329:full_adder port map (A => resultFA225, B => resultFA226, Cin => resultFA227, S => resultFA329, Cout => carryOutFA329);
FA330:full_adder port map (A => carryOutFA225, B => carryOutFA226, Cin => carryOutFA227, S => resultFA330, Cout => carryOutFA330);
FA331:full_adder port map (A => resultFA228, B => resultFA229, Cin => resultFA230, S => resultFA331, Cout => carryOutFA331);
FA332:full_adder port map (A => carryOutFA228, B => carryOutFA229, Cin => carryOutFA230, S => resultFA332, Cout => carryOutFA332);
FA333:full_adder port map (A => resultFA231, B => resultFA232, Cin => resultFA233, S => resultFA333, Cout => carryOutFA333);
FA334:full_adder port map (A => carryOutFA231, B => carryOutFA232, Cin => carryOutFA233, S => resultFA334, Cout => carryOutFA334);
FA335:full_adder port map (A => resultFA234, B => resultFA235, Cin => resultFA236, S => resultFA335, Cout => carryOutFA335);
FA336:full_adder port map (A => carryOutFA234, B => carryOutFA235, Cin => carryOutFA236, S => resultFA336, Cout => carryOutFA336);
FA337:full_adder port map (A => resultFA237, B => resultFA238, Cin => resultFA239, S => resultFA337, Cout => carryOutFA337);
FA338:full_adder port map (A => carryOutFA237, B => carryOutFA238, Cin => carryOutFA239, S => resultFA338, Cout => carryOutFA338);
FA339:full_adder port map (A => resultFA240, B => resultFA241, Cin => resultFA242, S => resultFA339, Cout => carryOutFA339);
FA340:full_adder port map (A => carryOutFA240, B => carryOutFA241, Cin => carryOutFA242, S => resultFA340, Cout => carryOutFA340);
FA341:full_adder port map (A => resultFA243, B => resultFA244, Cin => resultFA245, S => resultFA341, Cout => carryOutFA341);
FA342:full_adder port map (A => carryOutFA243, B => carryOutFA244, Cin => carryOutFA245, S => resultFA342, Cout => carryOutFA342);
FA343:full_adder port map (A => resultFA246, B => resultFA247, Cin => resultFA248, S => resultFA343, Cout => carryOutFA343);
FA344:full_adder port map (A => carryOutFA246, B => carryOutFA247, Cin => carryOutFA248, S => resultFA344, Cout => carryOutFA344);
FA345:full_adder port map (A => resultFA249, B => resultFA250, Cin => resultFA251, S => resultFA345, Cout => carryOutFA345);
FA346:full_adder port map (A => carryOutFA249, B => carryOutFA250, Cin => carryOutFA251, S => resultFA346, Cout => carryOutFA346);
FA347:full_adder port map (A => resultFA252, B => resultFA253, Cin => resultFA254, S => resultFA347, Cout => carryOutFA347);
FA348:full_adder port map (A => carryOutFA252, B => carryOutFA253, Cin => carryOutFA254, S => resultFA348, Cout => carryOutFA348);
FA349:full_adder port map (A => resultFA255, B => resultFA256, Cin => resultFA257, S => resultFA349, Cout => carryOutFA349);
FA350:full_adder port map (A => carryOutFA255, B => carryOutFA256, Cin => carryOutFA257, S => resultFA350, Cout => carryOutFA350);
FA351:full_adder port map (A => resultFA258, B => resultFA259, Cin => resultHA30, S => resultFA351, Cout => carryOutFA351);
FA352:full_adder port map (A => carryOutFA258, B => carryOutFA259, Cin => carryOutHA30, S => resultFA352, Cout => carryOutFA352);
FA353:full_adder port map (A => resultFA260, B => resultFA261, Cin => pp_ext(16)(23), S => resultFA353, Cout => carryOutFA353);
FA354:full_adder port map (A => carryOutFA260, B => carryOutFA261, Cin => resultFA262, S => resultFA354, Cout => carryOutFA354);
FA355:full_adder port map (A => resultHA31, B => pp_ext(15)(26), Cin => pp_ext(16)(24), S => resultFA355, Cout => carryOutFA355);
FA356:full_adder port map (A => carryOutFA262, B => carryOutHA31, Cin => resultFA263, S => resultFA356, Cout => carryOutFA356);
FA357:full_adder port map (A => pp_ext(14)(29), B => pp_ext(15)(27), Cin => pp_ext(16)(25), S => resultFA357, Cout => carryOutFA357);
FA358:full_adder port map (A => carryOutFA263, B => resultHA32, Cin => pp_ext(13)(32), S => resultFA358, Cout => carryOutFA358);
FA359:full_adder port map (A => pp_ext(14)(30), B => pp_ext(15)(28), Cin => pp_ext(16)(26), S => resultFA359, Cout => carryOutFA359);
FA360:full_adder port map (A => carryOutHA32, B => pp_ext(12)(35), Cin => pp_ext(13)(33), S => resultFA360, Cout => carryOutFA360);
FA361:full_adder port map (A => pp_ext(14)(31), B => pp_ext(15)(29), Cin => pp_ext(16)(27), S => resultFA361, Cout => carryOutFA361);
FA362:full_adder port map (A => pp_ext(12)(36), B => pp_ext(13)(34), Cin => pp_ext(14)(32), S => resultFA362, Cout => carryOutFA362);
HA37:half_adder port map (A => pp_ext(15)(30), B => pp_ext(16)(28), S => resultHA37, Cout => carryOutHA37);
FA363:full_adder port map (A => pp_ext(13)(35), B => pp_ext(14)(33), Cin => pp_ext(15)(31), S => resultFA363, Cout => carryOutFA363);
HA38:half_adder port map (A => pp_ext(13)(36), B => pp_ext(14)(34), S => resultHA38, Cout => carryOutHA38);
HA39:half_adder port map (A => pp_ext(0)(4), B => pp_ext(1)(4), S => resultHA39, Cout => carryOutHA39);
HA40:half_adder port map (A => pp_ext(0)(5), B => pp_ext(1)(5), S => resultHA40, Cout => carryOutHA40);
FA364:full_adder port map (A => resultHA33, B => pp_ext(2)(4), Cin => pp_ext(3)(2), S => resultFA364, Cout => carryOutFA364);
FA365:full_adder port map (A => carryOutHA33, B => resultHA34, Cin => pp_ext(2)(5), S => resultFA365, Cout => carryOutFA365);
FA366:full_adder port map (A => carryOutHA34, B => resultFA264, Cin => resultHA35, S => resultFA366, Cout => carryOutFA366);
FA367:full_adder port map (A => carryOutFA264, B => carryOutHA35, Cin => resultFA265, S => resultFA367, Cout => carryOutFA367);
FA368:full_adder port map (A => carryOutFA265, B => carryOutHA36, Cin => resultFA266, S => resultFA368, Cout => carryOutFA368);
FA369:full_adder port map (A => carryOutFA266, B => carryOutFA267, Cin => resultFA268, S => resultFA369, Cout => carryOutFA369);
FA370:full_adder port map (A => carryOutFA268, B => carryOutFA269, Cin => resultFA270, S => resultFA370, Cout => carryOutFA370);
FA371:full_adder port map (A => carryOutFA270, B => carryOutFA271, Cin => resultFA272, S => resultFA371, Cout => carryOutFA371);
FA372:full_adder port map (A => carryOutFA272, B => carryOutFA273, Cin => resultFA274, S => resultFA372, Cout => carryOutFA372);
FA373:full_adder port map (A => carryOutFA274, B => carryOutFA275, Cin => resultFA276, S => resultFA373, Cout => carryOutFA373);
FA374:full_adder port map (A => carryOutFA276, B => carryOutFA277, Cin => resultFA278, S => resultFA374, Cout => carryOutFA374);
FA375:full_adder port map (A => carryOutFA278, B => carryOutFA279, Cin => resultFA280, S => resultFA375, Cout => carryOutFA375);
FA376:full_adder port map (A => carryOutFA280, B => carryOutFA281, Cin => resultFA282, S => resultFA376, Cout => carryOutFA376);
FA377:full_adder port map (A => carryOutFA282, B => carryOutFA283, Cin => resultFA284, S => resultFA377, Cout => carryOutFA377);
FA378:full_adder port map (A => carryOutFA284, B => carryOutFA285, Cin => resultFA286, S => resultFA378, Cout => carryOutFA378);
FA379:full_adder port map (A => carryOutFA286, B => carryOutFA287, Cin => resultFA288, S => resultFA379, Cout => carryOutFA379);
FA380:full_adder port map (A => carryOutFA288, B => carryOutFA289, Cin => resultFA290, S => resultFA380, Cout => carryOutFA380);
FA381:full_adder port map (A => carryOutFA290, B => carryOutFA291, Cin => resultFA292, S => resultFA381, Cout => carryOutFA381);
FA382:full_adder port map (A => carryOutFA292, B => carryOutFA293, Cin => resultFA294, S => resultFA382, Cout => carryOutFA382);
FA383:full_adder port map (A => carryOutFA294, B => carryOutFA295, Cin => resultFA296, S => resultFA383, Cout => carryOutFA383);
FA384:full_adder port map (A => carryOutFA296, B => carryOutFA297, Cin => resultFA298, S => resultFA384, Cout => carryOutFA384);
FA385:full_adder port map (A => carryOutFA298, B => carryOutFA299, Cin => resultFA300, S => resultFA385, Cout => carryOutFA385);
FA386:full_adder port map (A => carryOutFA300, B => carryOutFA301, Cin => resultFA302, S => resultFA386, Cout => carryOutFA386);
FA387:full_adder port map (A => carryOutFA302, B => carryOutFA303, Cin => resultFA304, S => resultFA387, Cout => carryOutFA387);
FA388:full_adder port map (A => carryOutFA304, B => carryOutFA305, Cin => resultFA306, S => resultFA388, Cout => carryOutFA388);
FA389:full_adder port map (A => carryOutFA306, B => carryOutFA307, Cin => resultFA308, S => resultFA389, Cout => carryOutFA389);
FA390:full_adder port map (A => carryOutFA308, B => carryOutFA309, Cin => resultFA310, S => resultFA390, Cout => carryOutFA390);
FA391:full_adder port map (A => carryOutFA310, B => carryOutFA311, Cin => resultFA312, S => resultFA391, Cout => carryOutFA391);
FA392:full_adder port map (A => carryOutFA312, B => carryOutFA313, Cin => resultFA314, S => resultFA392, Cout => carryOutFA392);
FA393:full_adder port map (A => carryOutFA314, B => carryOutFA315, Cin => resultFA316, S => resultFA393, Cout => carryOutFA393);
FA394:full_adder port map (A => carryOutFA316, B => carryOutFA317, Cin => resultFA318, S => resultFA394, Cout => carryOutFA394);
FA395:full_adder port map (A => carryOutFA318, B => carryOutFA319, Cin => resultFA320, S => resultFA395, Cout => carryOutFA395);
FA396:full_adder port map (A => carryOutFA320, B => carryOutFA321, Cin => resultFA322, S => resultFA396, Cout => carryOutFA396);
FA397:full_adder port map (A => carryOutFA322, B => carryOutFA323, Cin => resultFA324, S => resultFA397, Cout => carryOutFA397);
FA398:full_adder port map (A => carryOutFA324, B => carryOutFA325, Cin => resultFA326, S => resultFA398, Cout => carryOutFA398);
FA399:full_adder port map (A => carryOutFA326, B => carryOutFA327, Cin => resultFA328, S => resultFA399, Cout => carryOutFA399);
FA400:full_adder port map (A => carryOutFA328, B => carryOutFA329, Cin => resultFA330, S => resultFA400, Cout => carryOutFA400);
FA401:full_adder port map (A => carryOutFA330, B => carryOutFA331, Cin => resultFA332, S => resultFA401, Cout => carryOutFA401);
FA402:full_adder port map (A => carryOutFA332, B => carryOutFA333, Cin => resultFA334, S => resultFA402, Cout => carryOutFA402);
FA403:full_adder port map (A => carryOutFA334, B => carryOutFA335, Cin => resultFA336, S => resultFA403, Cout => carryOutFA403);
FA404:full_adder port map (A => carryOutFA336, B => carryOutFA337, Cin => resultFA338, S => resultFA404, Cout => carryOutFA404);
FA405:full_adder port map (A => carryOutFA338, B => carryOutFA339, Cin => resultFA340, S => resultFA405, Cout => carryOutFA405);
FA406:full_adder port map (A => carryOutFA340, B => carryOutFA341, Cin => resultFA342, S => resultFA406, Cout => carryOutFA406);
FA407:full_adder port map (A => carryOutFA342, B => carryOutFA343, Cin => resultFA344, S => resultFA407, Cout => carryOutFA407);
FA408:full_adder port map (A => carryOutFA344, B => carryOutFA345, Cin => resultFA346, S => resultFA408, Cout => carryOutFA408);
FA409:full_adder port map (A => carryOutFA346, B => carryOutFA347, Cin => resultFA348, S => resultFA409, Cout => carryOutFA409);
FA410:full_adder port map (A => carryOutFA348, B => carryOutFA349, Cin => resultFA350, S => resultFA410, Cout => carryOutFA410);
FA411:full_adder port map (A => carryOutFA350, B => carryOutFA351, Cin => resultFA352, S => resultFA411, Cout => carryOutFA411);
FA412:full_adder port map (A => carryOutFA352, B => carryOutFA353, Cin => resultFA354, S => resultFA412, Cout => carryOutFA412);
FA413:full_adder port map (A => carryOutFA354, B => carryOutFA355, Cin => resultFA356, S => resultFA413, Cout => carryOutFA413);
FA414:full_adder port map (A => carryOutFA356, B => carryOutFA357, Cin => resultFA358, S => resultFA414, Cout => carryOutFA414);
FA415:full_adder port map (A => carryOutFA358, B => carryOutFA359, Cin => resultFA360, S => resultFA415, Cout => carryOutFA415);
FA416:full_adder port map (A => carryOutFA360, B => carryOutFA361, Cin => resultFA362, S => resultFA416, Cout => carryOutFA416);
FA417:full_adder port map (A => carryOutFA362, B => carryOutHA37, Cin => resultFA363, S => resultFA417, Cout => carryOutFA417);
FA418:full_adder port map (A => carryOutFA363, B => resultHA38, Cin => pp_ext(15)(32), S => resultFA418, Cout => carryOutFA418);
FA419:full_adder port map (A => carryOutHA38, B => pp_ext(14)(35), Cin => pp_ext(15)(33), S => resultFA419, Cout => carryOutFA419);
HA41:half_adder port map (A => pp_ext(14)(36), B => pp_ext(15)(34), S => resultHA41, Cout => carryOutHA41);
HA42:half_adder port map (A => pp_ext(0)(2), B => pp_ext(1)(2), S => resultHA42, Cout => carryOutHA42);
HA43:half_adder port map (A => pp_ext(0)(3), B => pp_ext(1)(3), S => resultHA43, Cout => carryOutHA43);
FA420:full_adder port map (A => resultHA39, B => pp_ext(2)(2), Cin => pp_ext(3)(0), S => resultFA420, Cout => carryOutFA420);
FA421:full_adder port map (A => carryOutHA39, B => resultHA40, Cin => pp_ext(2)(3), S => resultFA421, Cout => carryOutFA421);
FA422:full_adder port map (A => carryOutHA40, B => resultFA364, Cin => pp_ext(4)(0), S => resultFA422, Cout => carryOutFA422);
FA423:full_adder port map (A => carryOutFA364, B => resultFA365, Cin => pp_ext(3)(3), S => resultFA423, Cout => carryOutFA423);
FA424:full_adder port map (A => carryOutFA365, B => resultFA366, Cin => pp_ext(5)(0), S => resultFA424, Cout => carryOutFA424);
FA425:full_adder port map (A => carryOutFA366, B => resultFA367, Cin => resultHA36, S => resultFA425, Cout => carryOutFA425);
FA426:full_adder port map (A => carryOutFA367, B => resultFA368, Cin => resultFA267, S => resultFA426, Cout => carryOutFA426);
FA427:full_adder port map (A => carryOutFA368, B => resultFA369, Cin => resultFA269, S => resultFA427, Cout => carryOutFA427);
FA428:full_adder port map (A => carryOutFA369, B => resultFA370, Cin => resultFA271, S => resultFA428, Cout => carryOutFA428);
FA429:full_adder port map (A => carryOutFA370, B => resultFA371, Cin => resultFA273, S => resultFA429, Cout => carryOutFA429);
FA430:full_adder port map (A => carryOutFA371, B => resultFA372, Cin => resultFA275, S => resultFA430, Cout => carryOutFA430);
FA431:full_adder port map (A => carryOutFA372, B => resultFA373, Cin => resultFA277, S => resultFA431, Cout => carryOutFA431);
FA432:full_adder port map (A => carryOutFA373, B => resultFA374, Cin => resultFA279, S => resultFA432, Cout => carryOutFA432);
FA433:full_adder port map (A => carryOutFA374, B => resultFA375, Cin => resultFA281, S => resultFA433, Cout => carryOutFA433);
FA434:full_adder port map (A => carryOutFA375, B => resultFA376, Cin => resultFA283, S => resultFA434, Cout => carryOutFA434);
FA435:full_adder port map (A => carryOutFA376, B => resultFA377, Cin => resultFA285, S => resultFA435, Cout => carryOutFA435);
FA436:full_adder port map (A => carryOutFA377, B => resultFA378, Cin => resultFA287, S => resultFA436, Cout => carryOutFA436);
FA437:full_adder port map (A => carryOutFA378, B => resultFA379, Cin => resultFA289, S => resultFA437, Cout => carryOutFA437);
FA438:full_adder port map (A => carryOutFA379, B => resultFA380, Cin => resultFA291, S => resultFA438, Cout => carryOutFA438);
FA439:full_adder port map (A => carryOutFA380, B => resultFA381, Cin => resultFA293, S => resultFA439, Cout => carryOutFA439);
FA440:full_adder port map (A => carryOutFA381, B => resultFA382, Cin => resultFA295, S => resultFA440, Cout => carryOutFA440);
FA441:full_adder port map (A => carryOutFA382, B => resultFA383, Cin => resultFA297, S => resultFA441, Cout => carryOutFA441);
FA442:full_adder port map (A => carryOutFA383, B => resultFA384, Cin => resultFA299, S => resultFA442, Cout => carryOutFA442);
FA443:full_adder port map (A => carryOutFA384, B => resultFA385, Cin => resultFA301, S => resultFA443, Cout => carryOutFA443);
FA444:full_adder port map (A => carryOutFA385, B => resultFA386, Cin => resultFA303, S => resultFA444, Cout => carryOutFA444);
FA445:full_adder port map (A => carryOutFA386, B => resultFA387, Cin => resultFA305, S => resultFA445, Cout => carryOutFA445);
FA446:full_adder port map (A => carryOutFA387, B => resultFA388, Cin => resultFA307, S => resultFA446, Cout => carryOutFA446);
FA447:full_adder port map (A => carryOutFA388, B => resultFA389, Cin => resultFA309, S => resultFA447, Cout => carryOutFA447);
FA448:full_adder port map (A => carryOutFA389, B => resultFA390, Cin => resultFA311, S => resultFA448, Cout => carryOutFA448);
FA449:full_adder port map (A => carryOutFA390, B => resultFA391, Cin => resultFA313, S => resultFA449, Cout => carryOutFA449);
FA450:full_adder port map (A => carryOutFA391, B => resultFA392, Cin => resultFA315, S => resultFA450, Cout => carryOutFA450);
FA451:full_adder port map (A => carryOutFA392, B => resultFA393, Cin => resultFA317, S => resultFA451, Cout => carryOutFA451);
FA452:full_adder port map (A => carryOutFA393, B => resultFA394, Cin => resultFA319, S => resultFA452, Cout => carryOutFA452);
FA453:full_adder port map (A => carryOutFA394, B => resultFA395, Cin => resultFA321, S => resultFA453, Cout => carryOutFA453);
FA454:full_adder port map (A => carryOutFA395, B => resultFA396, Cin => resultFA323, S => resultFA454, Cout => carryOutFA454);
FA455:full_adder port map (A => carryOutFA396, B => resultFA397, Cin => resultFA325, S => resultFA455, Cout => carryOutFA455);
FA456:full_adder port map (A => carryOutFA397, B => resultFA398, Cin => resultFA327, S => resultFA456, Cout => carryOutFA456);
FA457:full_adder port map (A => carryOutFA398, B => resultFA399, Cin => resultFA329, S => resultFA457, Cout => carryOutFA457);
FA458:full_adder port map (A => carryOutFA399, B => resultFA400, Cin => resultFA331, S => resultFA458, Cout => carryOutFA458);
FA459:full_adder port map (A => carryOutFA400, B => resultFA401, Cin => resultFA333, S => resultFA459, Cout => carryOutFA459);
FA460:full_adder port map (A => carryOutFA401, B => resultFA402, Cin => resultFA335, S => resultFA460, Cout => carryOutFA460);
FA461:full_adder port map (A => carryOutFA402, B => resultFA403, Cin => resultFA337, S => resultFA461, Cout => carryOutFA461);
FA462:full_adder port map (A => carryOutFA403, B => resultFA404, Cin => resultFA339, S => resultFA462, Cout => carryOutFA462);
FA463:full_adder port map (A => carryOutFA404, B => resultFA405, Cin => resultFA341, S => resultFA463, Cout => carryOutFA463);
FA464:full_adder port map (A => carryOutFA405, B => resultFA406, Cin => resultFA343, S => resultFA464, Cout => carryOutFA464);
FA465:full_adder port map (A => carryOutFA406, B => resultFA407, Cin => resultFA345, S => resultFA465, Cout => carryOutFA465);
FA466:full_adder port map (A => carryOutFA407, B => resultFA408, Cin => resultFA347, S => resultFA466, Cout => carryOutFA466);
FA467:full_adder port map (A => carryOutFA408, B => resultFA409, Cin => resultFA349, S => resultFA467, Cout => carryOutFA467);
FA468:full_adder port map (A => carryOutFA409, B => resultFA410, Cin => resultFA351, S => resultFA468, Cout => carryOutFA468);
FA469:full_adder port map (A => carryOutFA410, B => resultFA411, Cin => resultFA353, S => resultFA469, Cout => carryOutFA469);
FA470:full_adder port map (A => carryOutFA411, B => resultFA412, Cin => resultFA355, S => resultFA470, Cout => carryOutFA470);
FA471:full_adder port map (A => carryOutFA412, B => resultFA413, Cin => resultFA357, S => resultFA471, Cout => carryOutFA471);
FA472:full_adder port map (A => carryOutFA413, B => resultFA414, Cin => resultFA359, S => resultFA472, Cout => carryOutFA472);
FA473:full_adder port map (A => carryOutFA414, B => resultFA415, Cin => resultFA361, S => resultFA473, Cout => carryOutFA473);
FA474:full_adder port map (A => carryOutFA415, B => resultFA416, Cin => resultHA37, S => resultFA474, Cout => carryOutFA474);
FA475:full_adder port map (A => carryOutFA416, B => resultFA417, Cin => pp_ext(16)(29), S => resultFA475, Cout => carryOutFA475);
FA476:full_adder port map (A => carryOutFA417, B => resultFA418, Cin => pp_ext(16)(30), S => resultFA476, Cout => carryOutFA476);
FA477:full_adder port map (A => carryOutFA418, B => resultFA419, Cin => pp_ext(16)(31), S => resultFA477, Cout => carryOutFA477);
FA478:full_adder port map (A => carryOutFA419, B => resultHA41, Cin => pp_ext(16)(32), S => resultFA478, Cout => carryOutFA478);
FA479:full_adder port map (A => carryOutHA41, B => pp_ext(15)(35), Cin => pp_ext(16)(33), S => resultFA479, Cout => carryOutFA479);
Addend1(0) <= pp_ext(0)(0);
Addend1(1) <= pp_ext(0)(1);
Addend1(2) <= resultHA42;
Addend1(3) <= carryOutHA42;
Addend1(4) <= carryOutHA43;
Addend1(5) <= carryOutFA420;
Addend1(6) <= carryOutFA421;
Addend1(7) <= carryOutFA422;
Addend1(8) <= carryOutFA423;
Addend1(9) <= carryOutFA424;
Addend1(10) <= carryOutFA425;
Addend1(11) <= carryOutFA426;
Addend1(12) <= carryOutFA427;
Addend1(13) <= carryOutFA428;
Addend1(14) <= carryOutFA429;
Addend1(15) <= carryOutFA430;
Addend1(16) <= carryOutFA431;
Addend1(17) <= carryOutFA432;
Addend1(18) <= carryOutFA433;
Addend1(19) <= carryOutFA434;
Addend1(20) <= carryOutFA435;
Addend1(21) <= carryOutFA436;
Addend1(22) <= carryOutFA437;
Addend1(23) <= carryOutFA438;
Addend1(24) <= carryOutFA439;
Addend1(25) <= carryOutFA440;
Addend1(26) <= carryOutFA441;
Addend1(27) <= carryOutFA442;
Addend1(28) <= carryOutFA443;
Addend1(29) <= carryOutFA444;
Addend1(30) <= carryOutFA445;
Addend1(31) <= carryOutFA446;
Addend1(32) <= carryOutFA447;
Addend1(33) <= carryOutFA448;
Addend1(34) <= carryOutFA449;
Addend1(35) <= carryOutFA450;
Addend1(36) <= carryOutFA451;
Addend1(37) <= carryOutFA452;
Addend1(38) <= carryOutFA453;
Addend1(39) <= carryOutFA454;
Addend1(40) <= carryOutFA455;
Addend1(41) <= carryOutFA456;
Addend1(42) <= carryOutFA457;
Addend1(43) <= carryOutFA458;
Addend1(44) <= carryOutFA459;
Addend1(45) <= carryOutFA460;
Addend1(46) <= carryOutFA461;
Addend1(47) <= carryOutFA462;
Addend1(48) <= carryOutFA463;
Addend1(49) <= carryOutFA464;
Addend1(50) <= carryOutFA465;
Addend1(51) <= carryOutFA466;
Addend1(52) <= carryOutFA467;
Addend1(53) <= carryOutFA468;
Addend1(54) <= carryOutFA469;
Addend1(55) <= carryOutFA470;
Addend1(56) <= carryOutFA471;
Addend1(57) <= carryOutFA472;
Addend1(58) <= carryOutFA473;
Addend1(59) <= carryOutFA474;
Addend1(60) <= carryOutFA475;
Addend1(61) <= carryOutFA476;
Addend1(62) <= carryOutFA477;
Addend1(63) <= carryOutFA478;
Addend2(0) <=pp_ext(1)(0);
Addend2(1) <= '0';
Addend2(2) <=pp_ext(2)(0);
Addend2(3) <=resultHA43;
Addend2(4) <=resultFA420;
Addend2(5) <=resultFA421;
Addend2(6) <=resultFA422;
Addend2(7) <=resultFA423;
Addend2(8) <=resultFA424;
Addend2(9) <=resultFA425;
Addend2(10) <=resultFA426;
Addend2(11) <=resultFA427;
Addend2(12) <=resultFA428;
Addend2(13) <=resultFA429;
Addend2(14) <=resultFA430;
Addend2(15) <=resultFA431;
Addend2(16) <=resultFA432;
Addend2(17) <=resultFA433;
Addend2(18) <=resultFA434;
Addend2(19) <=resultFA435;
Addend2(20) <=resultFA436;
Addend2(21) <=resultFA437;
Addend2(22) <=resultFA438;
Addend2(23) <=resultFA439;
Addend2(24) <=resultFA440;
Addend2(25) <=resultFA441;
Addend2(26) <=resultFA442;
Addend2(27) <=resultFA443;
Addend2(28) <=resultFA444;
Addend2(29) <=resultFA445;
Addend2(30) <=resultFA446;
Addend2(31) <=resultFA447;
Addend2(32) <=resultFA448;
Addend2(33) <=resultFA449;
Addend2(34) <=resultFA450;
Addend2(35) <=resultFA451;
Addend2(36) <=resultFA452;
Addend2(37) <=resultFA453;
Addend2(38) <=resultFA454;
Addend2(39) <=resultFA455;
Addend2(40) <=resultFA456;
Addend2(41) <=resultFA457;
Addend2(42) <=resultFA458;
Addend2(43) <=resultFA459;
Addend2(44) <=resultFA460;
Addend2(45) <=resultFA461;
Addend2(46) <=resultFA462;
Addend2(47) <=resultFA463;
Addend2(48) <=resultFA464;
Addend2(49) <=resultFA465;
Addend2(50) <=resultFA466;
Addend2(51) <=resultFA467;
Addend2(52) <=resultFA468;
Addend2(53) <=resultFA469;
Addend2(54) <=resultFA470;
Addend2(55) <=resultFA471;
Addend2(56) <=resultFA472;
Addend2(57) <=resultFA473;
Addend2(58) <=resultFA474;
Addend2(59) <=resultFA475;
Addend2(60) <=resultFA476;
Addend2(61) <=resultFA477;
Addend2(62) <=resultFA478;
Addend2(63) <=resultFA479;
end architecture;